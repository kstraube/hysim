library verilog;
use verilog.vl_types.all;
entity libio is
end libio;
