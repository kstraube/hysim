library verilog;
use verilog.vl_types.all;
entity libucode is
end libucode;
