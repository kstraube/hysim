library verilog;
use verilog.vl_types.all;
entity eth_tx_sv_unit is
end eth_tx_sv_unit;
