library verilog;
use verilog.vl_types.all;
entity exception_dma_sv_unit is
end exception_dma_sv_unit;
