library verilog;
use verilog.vl_types.all;
entity eth_rx_sv_unit is
end eth_rx_sv_unit;
