library verilog;
use verilog.vl_types.all;
entity itlbram_sv_unit is
end itlbram_sv_unit;
