library verilog;
use verilog.vl_types.all;
entity regacc_dma_sv_unit is
end regacc_dma_sv_unit;
