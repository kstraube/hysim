library verilog;
use verilog.vl_types.all;
entity libperfctr is
end libperfctr;
