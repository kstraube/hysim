library verilog;
use verilog.vl_types.all;
entity libxalu is
end libxalu;
