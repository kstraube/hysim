library verilog;
use verilog.vl_types.all;
entity dma_control_sv_unit is
end dma_control_sv_unit;
