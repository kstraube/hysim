library verilog;
use verilog.vl_types.all;
entity libconf is
end libconf;
