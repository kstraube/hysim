library verilog;
use verilog.vl_types.all;
entity pcie_blk_ll_tx is
    generic(
        TX_CPL_STALL_THRESHOLD: integer := 6;
        TX_DATACREDIT_FIX_EN: integer := 1;
        TX_DATACREDIT_FIX_1DWONLY: integer := 1;
        TX_DATACREDIT_FIX_MARGIN: integer := 6;
        MPS             : integer := 0;
        LEGACY_EP       : integer := 0
    );
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        trn_lnk_up_n    : in     vl_logic;
        llk_tx_data     : out    vl_logic_vector(63 downto 0);
        llk_tx_src_rdy_n: out    vl_logic;
        llk_tx_src_dsc_n: out    vl_logic;
        llk_tx_sof_n    : out    vl_logic;
        llk_tx_eof_n    : out    vl_logic;
        llk_tx_sop_n    : out    vl_logic;
        llk_tx_eop_n    : out    vl_logic;
        llk_tx_enable_n : out    vl_logic_vector(1 downto 0);
        llk_tx_ch_tc    : out    vl_logic_vector(2 downto 0);
        llk_tx_ch_fifo  : out    vl_logic_vector(1 downto 0);
        llk_tx_dst_rdy_n: in     vl_logic;
        llk_tx_chan_space: in     vl_logic_vector(9 downto 0);
        llk_tx_ch_posted_ready_n: in     vl_logic_vector(7 downto 0);
        llk_tx_ch_non_posted_ready_n: in     vl_logic_vector(7 downto 0);
        llk_tx_ch_completion_ready_n: in     vl_logic_vector(7 downto 0);
        trn_td          : in     vl_logic_vector(63 downto 0);
        trn_trem_n      : in     vl_logic_vector(7 downto 0);
        trn_tsof_n      : in     vl_logic;
        trn_teof_n      : in     vl_logic;
        trn_tsrc_rdy_n  : in     vl_logic;
        trn_tsrc_dsc_n  : in     vl_logic;
        trn_terrfwd_n   : in     vl_logic;
        trn_tdst_rdy_n  : out    vl_logic;
        trn_tdst_dsc_n  : out    vl_logic;
        trn_tbuf_av_cpl : out    vl_logic;
        tx_ch_credits_consumed: in     vl_logic_vector(7 downto 0);
        tx_pd_credits_available: in     vl_logic_vector(11 downto 0);
        tx_pd_credits_consumed: in     vl_logic_vector(11 downto 0);
        tx_npd_credits_available: in     vl_logic_vector(11 downto 0);
        tx_npd_credits_consumed: in     vl_logic_vector(11 downto 0);
        tx_cd_credits_available: in     vl_logic_vector(11 downto 0);
        tx_cd_credits_consumed: in     vl_logic_vector(11 downto 0);
        clear_cpl_count : out    vl_logic;
        pd_credit_limited: in     vl_logic;
        npd_credit_limited: in     vl_logic;
        cd_credit_limited: in     vl_logic;
        trn_pfc_cplh_cl_upd: in     vl_logic;
        trn_pfc_cplh_cl : in     vl_logic_vector(7 downto 0);
        max_payload_size: in     vl_logic_vector(2 downto 0);
        l0_stats_cfg_transmitted: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of TX_CPL_STALL_THRESHOLD : constant is 1;
    attribute mti_svvh_generic_type of TX_DATACREDIT_FIX_EN : constant is 1;
    attribute mti_svvh_generic_type of TX_DATACREDIT_FIX_1DWONLY : constant is 1;
    attribute mti_svvh_generic_type of TX_DATACREDIT_FIX_MARGIN : constant is 1;
    attribute mti_svvh_generic_type of MPS : constant is 1;
    attribute mti_svvh_generic_type of LEGACY_EP : constant is 1;
end pcie_blk_ll_tx;
