library verilog;
use verilog.vl_types.all;
entity immu_sv_unit is
end immu_sv_unit;
