library verilog;
use verilog.vl_types.all;
entity libmemif_sv_unit is
end libmemif_sv_unit;
