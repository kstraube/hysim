library verilog;
use verilog.vl_types.all;
entity icache_sv_unit is
end icache_sv_unit;
