library verilog;
use verilog.vl_types.all;
entity microcode_sv_unit is
end microcode_sv_unit;
