library verilog;
use verilog.vl_types.all;
entity libtm is
end libtm;
