library verilog;
use verilog.vl_types.all;
entity decode_sv_unit is
end decode_sv_unit;
