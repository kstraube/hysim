library verilog;
use verilog.vl_types.all;
entity libmmu_sv_unit is
end libmmu_sv_unit;
