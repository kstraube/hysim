library verilog;
use verilog.vl_types.all;
entity udcache_nb_mmu_sv_unit is
end udcache_nb_mmu_sv_unit;
