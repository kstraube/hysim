library verilog;
use verilog.vl_types.all;
entity mac_fedriver_sv_unit is
end mac_fedriver_sv_unit;
