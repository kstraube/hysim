library verilog;
use verilog.vl_types.all;
entity pcie_blk_cf_mgmt is
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        completer_id    : in     vl_logic_vector(12 downto 0);
        mgmt_addr       : out    vl_logic_vector(10 downto 0);
        mgmt_wren       : out    vl_logic;
        mgmt_rden       : out    vl_logic;
        mgmt_wdata      : out    vl_logic_vector(31 downto 0);
        mgmt_bwren      : out    vl_logic_vector(3 downto 0);
        mgmt_rdata      : in     vl_logic_vector(31 downto 0);
        mgmt_pso        : in     vl_logic_vector(16 downto 0);
        cfg_dsn         : in     vl_logic_vector(63 downto 0);
        cfg_do          : out    vl_logic_vector(31 downto 0);
        cfg_rd_wr_done_n: out    vl_logic;
        cfg_dwaddr      : in     vl_logic_vector(11 downto 0);
        cfg_rd_en_n     : in     vl_logic;
        cfg_rx_bar0     : out    vl_logic_vector(31 downto 0);
        cfg_rx_bar1     : out    vl_logic_vector(31 downto 0);
        cfg_rx_bar2     : out    vl_logic_vector(31 downto 0);
        cfg_rx_bar3     : out    vl_logic_vector(31 downto 0);
        cfg_rx_bar4     : out    vl_logic_vector(31 downto 0);
        cfg_rx_bar5     : out    vl_logic_vector(31 downto 0);
        cfg_rx_xrom     : out    vl_logic_vector(31 downto 0);
        cfg_status      : out    vl_logic_vector(15 downto 0);
        cfg_command     : out    vl_logic_vector(15 downto 0);
        cfg_dstatus     : out    vl_logic_vector(15 downto 0);
        cfg_dcommand    : out    vl_logic_vector(15 downto 0);
        cfg_lstatus     : out    vl_logic_vector(15 downto 0);
        cfg_lcommand    : out    vl_logic_vector(15 downto 0);
        cfg_pmcsr       : out    vl_logic_vector(31 downto 0);
        cfg_dcap        : out    vl_logic_vector(31 downto 0);
        cfg_msgctrl     : out    vl_logic_vector(15 downto 0);
        cfg_msgladdr    : out    vl_logic_vector(31 downto 0);
        cfg_msguaddr    : out    vl_logic_vector(31 downto 0);
        cfg_msgdata     : out    vl_logic_vector(15 downto 0);
        cfg_bus_number  : out    vl_logic_vector(7 downto 0);
        cfg_device_number: out    vl_logic_vector(4 downto 0);
        cfg_function_number: out    vl_logic_vector(2 downto 0);
        llk_rx_data_d   : in     vl_logic_vector(63 downto 0);
        llk_rx_src_rdy_n: in     vl_logic;
        l0_dll_error_vector: in     vl_logic_vector(6 downto 0);
        l0_rx_mac_link_error: in     vl_logic_vector(1 downto 0);
        l0_stats_cfg_received: in     vl_logic;
        l0_stats_cfg_transmitted: in     vl_logic;
        l0_set_unsupported_request_other_error: in     vl_logic;
        l0_set_detected_corr_error: in     vl_logic
    );
end pcie_blk_cf_mgmt;
