library verilog;
use verilog.vl_types.all;
entity mt16htf25664hy_sv_unit is
end mt16htf25664hy_sv_unit;
