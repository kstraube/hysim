library verilog;
use verilog.vl_types.all;
entity perfctr_sv_unit is
end perfctr_sv_unit;
