library verilog;
use verilog.vl_types.all;
entity dtlbram_sv_unit is
end dtlbram_sv_unit;
