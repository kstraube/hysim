library verilog;
use verilog.vl_types.all;
entity eth_tm_control_sv_unit is
end eth_tm_control_sv_unit;
