library verilog;
use verilog.vl_types.all;
entity dtlb_2way_split_sv_unit is
end dtlb_2way_split_sv_unit;
