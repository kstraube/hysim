library verilog;
use verilog.vl_types.all;
entity top_1P_bee3_neweth_sv_unit is
end top_1P_bee3_neweth_sv_unit;
