library verilog;
use verilog.vl_types.all;
entity dramctrl_network_sv_unit is
end dramctrl_network_sv_unit;
