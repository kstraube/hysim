library verilog;
use verilog.vl_types.all;
entity xalu_fast_sv_unit is
end xalu_fast_sv_unit;
