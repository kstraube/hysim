library verilog;
use verilog.vl_types.all;
entity tm_cpu_l1_ring_sv_unit is
end tm_cpu_l1_ring_sv_unit;
