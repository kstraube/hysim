library verilog;
use verilog.vl_types.all;
entity pcie_blk_cf is
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        trn_lnk_up_n    : out    vl_logic;
        mac_link_up     : in     vl_logic;
        mac_negotiated_link_width: in     vl_logic_vector(3 downto 0);
        llk_tc_status   : in     vl_logic_vector(7 downto 0);
        io_space_enable : in     vl_logic;
        mem_space_enable: in     vl_logic;
        bus_master_enable: in     vl_logic;
        parity_error_response: in     vl_logic;
        serr_enable     : in     vl_logic;
        msi_enable      : in     vl_logic;
        completer_id    : in     vl_logic_vector(12 downto 0);
        max_read_request_size: in     vl_logic_vector(2 downto 0);
        max_payload_size: in     vl_logic_vector(2 downto 0);
        legacy_int_request: out    vl_logic;
        transactions_pending: out    vl_logic;
        msi_request     : out    vl_logic_vector(3 downto 0);
        cfg_interrupt_assert_n: in     vl_logic;
        cfg_interrupt_di: in     vl_logic_vector(7 downto 0);
        cfg_interrupt_mmenable: out    vl_logic_vector(2 downto 0);
        cfg_interrupt_msienable: out    vl_logic;
        cfg_interrupt_do: out    vl_logic_vector(7 downto 0);
        msi_8bit_en     : in     vl_logic;
        mgmt_addr       : out    vl_logic_vector(10 downto 0);
        mgmt_wren       : out    vl_logic;
        mgmt_rden       : out    vl_logic;
        mgmt_wdata      : out    vl_logic_vector(31 downto 0);
        mgmt_bwren      : out    vl_logic_vector(3 downto 0);
        mgmt_rdata      : in     vl_logic_vector(31 downto 0);
        mgmt_pso        : in     vl_logic_vector(16 downto 0);
        llk_rx_data_d   : in     vl_logic_vector(63 downto 0);
        llk_rx_src_rdy_n: in     vl_logic;
        l0_stats_cfg_received: in     vl_logic;
        l0_stats_cfg_transmitted: in     vl_logic;
        cfg_do          : out    vl_logic_vector(31 downto 0);
        cfg_di          : in     vl_logic_vector(31 downto 0);
        cfg_dsn         : in     vl_logic_vector(63 downto 0);
        cfg_byte_en_n   : in     vl_logic_vector(3 downto 0);
        cfg_dwaddr      : in     vl_logic_vector(11 downto 0);
        cfg_rd_wr_done_n: out    vl_logic;
        cfg_wr_en_n     : in     vl_logic;
        cfg_rd_en_n     : in     vl_logic;
        cfg_err_cor_n   : in     vl_logic;
        cfg_err_ur_n    : in     vl_logic;
        cfg_err_ecrc_n  : in     vl_logic;
        cfg_err_cpl_timeout_n: in     vl_logic;
        cfg_err_cpl_abort_n: in     vl_logic;
        cfg_err_cpl_unexpect_n: in     vl_logic;
        cfg_err_posted_n: in     vl_logic;
        cfg_err_locked_n: in     vl_logic;
        cfg_interrupt_n : in     vl_logic;
        cfg_interrupt_rdy_n: out    vl_logic;
        cfg_turnoff_ok_n: in     vl_logic;
        cfg_to_turnoff_n: out    vl_logic;
        cfg_pm_wake_n   : in     vl_logic;
        cfg_err_tlp_cpl_header: in     vl_logic_vector(47 downto 0);
        cfg_err_cpl_rdy_n: out    vl_logic;
        cfg_trn_pending_n: in     vl_logic;
        cfg_rx_bar0     : out    vl_logic_vector(31 downto 0);
        cfg_rx_bar1     : out    vl_logic_vector(31 downto 0);
        cfg_rx_bar2     : out    vl_logic_vector(31 downto 0);
        cfg_rx_bar3     : out    vl_logic_vector(31 downto 0);
        cfg_rx_bar4     : out    vl_logic_vector(31 downto 0);
        cfg_rx_bar5     : out    vl_logic_vector(31 downto 0);
        cfg_rx_xrom     : out    vl_logic_vector(31 downto 0);
        cfg_status      : out    vl_logic_vector(15 downto 0);
        cfg_command     : out    vl_logic_vector(15 downto 0);
        cfg_dstatus     : out    vl_logic_vector(15 downto 0);
        cfg_dcommand    : out    vl_logic_vector(15 downto 0);
        cfg_lstatus     : out    vl_logic_vector(15 downto 0);
        cfg_lcommand    : out    vl_logic_vector(15 downto 0);
        cfg_pmcsr       : out    vl_logic_vector(31 downto 0);
        cfg_dcap        : out    vl_logic_vector(31 downto 0);
        cfg_bus_number  : out    vl_logic_vector(7 downto 0);
        cfg_device_number: out    vl_logic_vector(4 downto 0);
        cfg_function_number: out    vl_logic_vector(2 downto 0);
        cfg_pcie_link_state_n: out    vl_logic_vector(2 downto 0);
        rx_err_cpl_ep_n : in     vl_logic;
        tx_err_wr_ep_n  : in     vl_logic;
        rx_err_ep_n     : in     vl_logic;
        rx_err_tlp_poisoned_n: in     vl_logic;
        rx_err_cpl_abort_n: in     vl_logic;
        rx_err_cpl_ur_n : in     vl_logic;
        rx_err_tlp_ur_n : in     vl_logic;
        rx_err_tlp_ur_lock_n: in     vl_logic;
        rx_err_tlp_p_cpl_n: in     vl_logic;
        rx_err_tlp_malformed_n: in     vl_logic;
        rx_err_tlp_hdr  : in     vl_logic_vector(47 downto 0);
        cfg_arb_td      : out    vl_logic_vector(63 downto 0);
        cfg_arb_trem_n  : out    vl_logic_vector(7 downto 0);
        cfg_arb_tsof_n  : out    vl_logic;
        cfg_arb_teof_n  : out    vl_logic;
        cfg_arb_tsrc_rdy_n: out    vl_logic;
        cfg_arb_tdst_rdy_n: in     vl_logic;
        l0_dll_error_vector: in     vl_logic_vector(6 downto 0);
        l0_rx_mac_link_error: in     vl_logic_vector(1 downto 0);
        l0_set_unsupported_request_other_error: out    vl_logic;
        l0_set_detected_fatal_error: out    vl_logic;
        l0_set_detected_nonfatal_error: out    vl_logic;
        l0_set_detected_corr_error: out    vl_logic;
        l0_set_user_system_error: out    vl_logic;
        l0_set_user_master_data_parity: out    vl_logic;
        l0_set_user_signaled_target_abort: out    vl_logic;
        l0_set_user_received_target_abort: out    vl_logic;
        l0_set_user_received_master_abort: out    vl_logic;
        l0_set_user_detected_parity_error: out    vl_logic;
        l0_ltssm_state  : in     vl_logic_vector(3 downto 0);
        l0_pwr_turn_off_req: in     vl_logic;
        l0_pme_req_in   : out    vl_logic;
        l0_pme_ack      : in     vl_logic
    );
end pcie_blk_cf;
