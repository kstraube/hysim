library verilog;
use verilog.vl_types.all;
entity fpu_sv_unit is
end fpu_sv_unit;
