library verilog;
use verilog.vl_types.all;
entity speed_tm_sv_unit is
end speed_tm_sv_unit;
