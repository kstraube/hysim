library verilog;
use verilog.vl_types.all;
entity ReadModule_sv_unit is
end ReadModule_sv_unit;
