library verilog;
use verilog.vl_types.all;
entity pcie_blk_cf_arb is
    generic(
        st_reset        : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        st_clear_count  : vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi0, Hi1);
        st_clear_send   : vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi1, Hi0);
        st_cleared_all  : vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi1, Hi1);
        st_cplu_req     : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        st_cplt_req     : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi0);
        st_ftl_req      : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi1);
        st_nfl_req      : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi0, Hi0);
        st_cor_req      : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi0, Hi1);
        st_send_pm      : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi1, Hi0);
        st_send_msi_32  : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi1, Hi1);
        st_send_msi_64  : vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi0, Hi0);
        st_code_send_asrt: vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi0, Hi0);
        st_code_send_d_asrt: vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi0, Hi1);
        type_msg_intr   : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi0, Hi0);
        UR              : vl_logic := Hi0;
        CA              : vl_logic := Hi1;
        LOCK            : vl_logic := Hi0;
        rsvd_BYTE0      : vl_logic := Hi0;
        fmt_mwr_3dwhdr_data: vl_logic_vector(0 to 1) := (Hi1, Hi0);
        fmt_mwr_4dwhdr_data: vl_logic_vector(0 to 1) := (Hi1, Hi1);
        fmt_msg         : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        fmt_cpl         : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        type_mwr        : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        type_msg        : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi0);
        type_cpl        : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi0);
        type_cpllock    : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi1);
        rsvd_msb_BYTE1  : vl_logic := Hi0;
        tc_param        : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        rsvd_BYTE1      : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        td              : vl_logic := Hi0;
        ep              : vl_logic := Hi0;
        attr_param      : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        rsvd_BYTE2      : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        len_98          : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        len_70_BYTE3    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        len_70_mwrd_BYTE3: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        compl_status_sc : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        compl_status_ur : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        compl_status_ca : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        bcm             : vl_logic := Hi0;
        msg_code_err_cor_BYTE7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        msg_code_err_nfl_BYTE7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1);
        msg_code_err_ftl_BYTE7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1);
        rsvd_BYTE11     : vl_logic := Hi0;
        msg_code_pm_pme_BYTE7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        msg_code_pme_to_ack_BYTE7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1);
        type_msg_pme_to_ack: vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi0, Hi1);
        last_dw_byte_enable_BYTE7: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        first_dw_byte_enable_BYTE7: vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        msg_code_asrt_inta_BYTE7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        msg_code_asrt_intb_BYTE7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        msg_code_asrt_intc_BYTE7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0);
        msg_code_asrt_intd_BYTE7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        msg_code_d_asrt_inta_BYTE7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        msg_code_d_asrt_intb_BYTE7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1);
        msg_code_d_asrt_intc_BYTE7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        msg_code_d_asrt_intd_BYTE7: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        TX_IDLE         : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        TX_DW1          : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        TX_DW3          : vl_logic_vector(0 to 1) := (Hi1, Hi0);
        SEND_GRANT      : vl_logic_vector(0 to 1) := (Hi1, Hi1)
    );
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        cfg_bus_number  : in     vl_logic_vector(7 downto 0);
        cfg_device_number: in     vl_logic_vector(4 downto 0);
        cfg_function_number: in     vl_logic_vector(2 downto 0);
        msi_data        : in     vl_logic_vector(15 downto 0);
        msi_laddr       : in     vl_logic_vector(31 downto 0);
        msi_haddr       : in     vl_logic_vector(31 downto 0);
        send_cor        : in     vl_logic;
        send_nfl        : in     vl_logic;
        send_ftl        : in     vl_logic;
        send_cplt       : in     vl_logic;
        send_cplu       : in     vl_logic;
        cmt_rd_hdr      : in     vl_logic_vector(49 downto 0);
        cfg_rd_hdr      : in     vl_logic_vector(49 downto 0);
        request_data    : out    vl_logic_vector(49 downto 0);
        grant           : out    vl_logic;
        cs_is_cplu      : out    vl_logic;
        cs_is_cplt      : out    vl_logic;
        cs_is_cor       : out    vl_logic;
        cs_is_nfl       : out    vl_logic;
        cs_is_ftl       : out    vl_logic;
        cs_is_pm        : out    vl_logic;
        send_pmeack     : in     vl_logic;
        cs_is_intr      : out    vl_logic;
        intr_vector     : in     vl_logic_vector(7 downto 0);
        intr_req_type   : in     vl_logic_vector(1 downto 0);
        intr_req_valid  : in     vl_logic;
        cfg_arb_td      : out    vl_logic_vector(63 downto 0);
        cfg_arb_trem_n  : out    vl_logic_vector(7 downto 0);
        cfg_arb_tsof_n  : out    vl_logic;
        cfg_arb_teof_n  : out    vl_logic;
        cfg_arb_tsrc_rdy_n: out    vl_logic;
        cfg_arb_tdst_rdy_n: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of st_reset : constant is 2;
    attribute mti_svvh_generic_type of st_clear_count : constant is 2;
    attribute mti_svvh_generic_type of st_clear_send : constant is 2;
    attribute mti_svvh_generic_type of st_cleared_all : constant is 2;
    attribute mti_svvh_generic_type of st_cplu_req : constant is 2;
    attribute mti_svvh_generic_type of st_cplt_req : constant is 2;
    attribute mti_svvh_generic_type of st_ftl_req : constant is 2;
    attribute mti_svvh_generic_type of st_nfl_req : constant is 2;
    attribute mti_svvh_generic_type of st_cor_req : constant is 2;
    attribute mti_svvh_generic_type of st_send_pm : constant is 2;
    attribute mti_svvh_generic_type of st_send_msi_32 : constant is 2;
    attribute mti_svvh_generic_type of st_send_msi_64 : constant is 2;
    attribute mti_svvh_generic_type of st_code_send_asrt : constant is 2;
    attribute mti_svvh_generic_type of st_code_send_d_asrt : constant is 2;
    attribute mti_svvh_generic_type of type_msg_intr : constant is 1;
    attribute mti_svvh_generic_type of UR : constant is 1;
    attribute mti_svvh_generic_type of CA : constant is 1;
    attribute mti_svvh_generic_type of LOCK : constant is 1;
    attribute mti_svvh_generic_type of rsvd_BYTE0 : constant is 1;
    attribute mti_svvh_generic_type of fmt_mwr_3dwhdr_data : constant is 1;
    attribute mti_svvh_generic_type of fmt_mwr_4dwhdr_data : constant is 1;
    attribute mti_svvh_generic_type of fmt_msg : constant is 1;
    attribute mti_svvh_generic_type of fmt_cpl : constant is 1;
    attribute mti_svvh_generic_type of type_mwr : constant is 1;
    attribute mti_svvh_generic_type of type_msg : constant is 1;
    attribute mti_svvh_generic_type of type_cpl : constant is 1;
    attribute mti_svvh_generic_type of type_cpllock : constant is 1;
    attribute mti_svvh_generic_type of rsvd_msb_BYTE1 : constant is 1;
    attribute mti_svvh_generic_type of tc_param : constant is 1;
    attribute mti_svvh_generic_type of rsvd_BYTE1 : constant is 1;
    attribute mti_svvh_generic_type of td : constant is 1;
    attribute mti_svvh_generic_type of ep : constant is 1;
    attribute mti_svvh_generic_type of attr_param : constant is 1;
    attribute mti_svvh_generic_type of rsvd_BYTE2 : constant is 1;
    attribute mti_svvh_generic_type of len_98 : constant is 1;
    attribute mti_svvh_generic_type of len_70_BYTE3 : constant is 1;
    attribute mti_svvh_generic_type of len_70_mwrd_BYTE3 : constant is 1;
    attribute mti_svvh_generic_type of compl_status_sc : constant is 1;
    attribute mti_svvh_generic_type of compl_status_ur : constant is 1;
    attribute mti_svvh_generic_type of compl_status_ca : constant is 1;
    attribute mti_svvh_generic_type of bcm : constant is 1;
    attribute mti_svvh_generic_type of msg_code_err_cor_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of msg_code_err_nfl_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of msg_code_err_ftl_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of rsvd_BYTE11 : constant is 1;
    attribute mti_svvh_generic_type of msg_code_pm_pme_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of msg_code_pme_to_ack_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of type_msg_pme_to_ack : constant is 1;
    attribute mti_svvh_generic_type of last_dw_byte_enable_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of first_dw_byte_enable_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of msg_code_asrt_inta_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of msg_code_asrt_intb_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of msg_code_asrt_intc_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of msg_code_asrt_intd_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of msg_code_d_asrt_inta_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of msg_code_d_asrt_intb_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of msg_code_d_asrt_intc_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of msg_code_d_asrt_intd_BYTE7 : constant is 1;
    attribute mti_svvh_generic_type of TX_IDLE : constant is 1;
    attribute mti_svvh_generic_type of TX_DW1 : constant is 1;
    attribute mti_svvh_generic_type of TX_DW3 : constant is 1;
    attribute mti_svvh_generic_type of SEND_GRANT : constant is 1;
end pcie_blk_cf_arb;
