library verilog;
use verilog.vl_types.all;
entity libtech is
end libtech;
