library verilog;
use verilog.vl_types.all;
entity tm_cache_sv_unit is
end tm_cache_sv_unit;
