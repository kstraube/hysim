library verilog;
use verilog.vl_types.all;
entity prod_fixes is
    generic(
        STATE_SIZE      : integer := 5;
        ALGN            : vl_logic_vector;
        Q_TS            : vl_logic_vector;
        SYM2            : vl_logic_vector;
        SYM3            : vl_logic_vector;
        SYM4            : vl_logic_vector;
        PAD             : vl_logic_vector(8 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1);
        COM             : vl_logic_vector(8 downto 0) := (Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        SKP             : vl_logic_vector(8 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        IDL             : vl_logic_vector(8 downto 0) := (Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        SDP             : vl_logic_vector(8 downto 0) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        \END\           : vl_logic_vector(8 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1);
        LT_POLLING      : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi0);
        LT_CONFIG       : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi1);
        LT_L0           : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi0, Hi0);
        LT_RECOVERY     : vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi0, Hi0);
        IS_D            : vl_logic := Hi0;
        IS_K            : vl_logic := Hi1
    );
    port(
        clk             : in     vl_logic;
        bit_reset_n     : in     vl_logic;
        l0_ltssm_state  : in     vl_logic_vector(3 downto 0);
        chan_bond_done  : in     vl_logic;
        negotiated_link_width: in     vl_logic_vector(3 downto 0);
        trn_lnk_up_n    : in     vl_logic;
        pipe_rx_data_k  : in     vl_logic_vector(7 downto 0);
        pipe_rx_valid   : in     vl_logic_vector(7 downto 0);
        pipe_rx_data_l0 : in     vl_logic_vector(7 downto 0);
        pipe_rx_data_l1 : in     vl_logic_vector(7 downto 0);
        pipe_rx_data_l2 : in     vl_logic_vector(7 downto 0);
        pipe_rx_data_l3 : in     vl_logic_vector(7 downto 0);
        pipe_rx_data_l4 : in     vl_logic_vector(7 downto 0);
        pipe_rx_data_l5 : in     vl_logic_vector(7 downto 0);
        pipe_rx_data_l6 : in     vl_logic_vector(7 downto 0);
        pipe_rx_data_l7 : in     vl_logic_vector(7 downto 0);
        pipe_rx_data_l0_out: out    vl_logic_vector(7 downto 0);
        pipe_rx_data_l1_out: out    vl_logic_vector(7 downto 0);
        pipe_rx_data_l2_out: out    vl_logic_vector(7 downto 0);
        pipe_rx_data_l3_out: out    vl_logic_vector(7 downto 0);
        pipe_rx_data_l4_out: out    vl_logic_vector(7 downto 0);
        pipe_rx_data_l5_out: out    vl_logic_vector(7 downto 0);
        pipe_rx_data_l6_out: out    vl_logic_vector(7 downto 0);
        pipe_rx_data_l7_out: out    vl_logic_vector(7 downto 0);
        upcfgcap_cycle  : out    vl_logic;
        masking_ack     : out    vl_logic;
        pipe_rx_data_k_out: out    vl_logic_vector(7 downto 0);
        pipe_rx_valid_out: out    vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of STATE_SIZE : constant is 1;
    attribute mti_svvh_generic_type of ALGN : constant is 4;
    attribute mti_svvh_generic_type of Q_TS : constant is 4;
    attribute mti_svvh_generic_type of SYM2 : constant is 4;
    attribute mti_svvh_generic_type of SYM3 : constant is 4;
    attribute mti_svvh_generic_type of SYM4 : constant is 4;
    attribute mti_svvh_generic_type of PAD : constant is 2;
    attribute mti_svvh_generic_type of COM : constant is 2;
    attribute mti_svvh_generic_type of SKP : constant is 2;
    attribute mti_svvh_generic_type of IDL : constant is 2;
    attribute mti_svvh_generic_type of SDP : constant is 2;
    attribute mti_svvh_generic_type of \END\ : constant is 2;
    attribute mti_svvh_generic_type of LT_POLLING : constant is 2;
    attribute mti_svvh_generic_type of LT_CONFIG : constant is 2;
    attribute mti_svvh_generic_type of LT_L0 : constant is 2;
    attribute mti_svvh_generic_type of LT_RECOVERY : constant is 2;
    attribute mti_svvh_generic_type of IS_D : constant is 1;
    attribute mti_svvh_generic_type of IS_K : constant is 1;
end prod_fixes;
