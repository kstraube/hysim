library verilog;
use verilog.vl_types.all;
entity debugdma_sv_unit is
end debugdma_sv_unit;
