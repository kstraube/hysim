library verilog;
use verilog.vl_types.all;
entity WriteModule2_sv_unit is
end WriteModule2_sv_unit;
