library verilog;
use verilog.vl_types.all;
entity irqmp_sv_unit is
end irqmp_sv_unit;
