library verilog;
use verilog.vl_types.all;
entity libcache is
end libcache;
