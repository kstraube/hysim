library verilog;
use verilog.vl_types.all;
entity tm_cpu_dram_gsf_sv_unit is
end tm_cpu_dram_gsf_sv_unit;
