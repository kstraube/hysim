library verilog;
use verilog.vl_types.all;
entity alulogic_sv_unit is
end alulogic_sv_unit;
