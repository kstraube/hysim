library verilog;
use verilog.vl_types.all;
entity fpregfile_sv_unit is
end fpregfile_sv_unit;
