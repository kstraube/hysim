library verilog;
use verilog.vl_types.all;
entity ifetch_dma_sv_unit is
end ifetch_dma_sv_unit;
