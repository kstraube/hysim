library verilog;
use verilog.vl_types.all;
entity tlm_rx_data_snk is
    generic(
        DW              : integer := 32;
        FCW             : integer := 6;
        BARW            : integer := 7;
        DOWNSTREAM_PORT : integer := 0;
        MPS             : integer := 512;
        TYPE1_UR        : integer := 0
    );
    port(
        clk_i           : in     vl_logic;
        reset_i         : in     vl_logic;
        d_o             : out    vl_logic_vector;
        sof_o           : out    vl_logic;
        eof_o           : out    vl_logic;
        preeof_o        : out    vl_logic;
        src_rdy_o       : out    vl_logic;
        rem_o           : out    vl_logic;
        dsc_o           : out    vl_logic;
        cfg_o           : out    vl_logic;
        np_o            : out    vl_logic;
        cpl_o           : out    vl_logic;
        locked_o        : out    vl_logic;
        bar_o           : out    vl_logic_vector;
        rid_o           : out    vl_logic;
        vend_msg_o      : out    vl_logic;
        bar_src_rdy_o   : out    vl_logic;
        fc_use_p_o      : out    vl_logic;
        fc_use_np_o     : out    vl_logic;
        fc_use_cpl_o    : out    vl_logic;
        fc_use_data_o   : out    vl_logic_vector;
        fc_unuse_o      : out    vl_logic;
        d_i             : in     vl_logic_vector;
        sof_i           : in     vl_logic;
        eof_i           : in     vl_logic;
        rem_i           : in     vl_logic;
        src_rdy_i       : in     vl_logic;
        src_dsc_i       : in     vl_logic;
        vc_hit_o        : out    vl_logic;
        pm_as_nak_l1_o  : out    vl_logic;
        pm_turn_off_o   : out    vl_logic;
        pm_set_slot_pwr_o: out    vl_logic;
        pm_set_slot_pwr_data_o: out    vl_logic_vector(9 downto 0);
        pm_suspend_req_i: in     vl_logic;
        err_tlp_cpl_header_o: out    vl_logic_vector(47 downto 0);
        err_tlp_p_o     : out    vl_logic;
        err_tlp_ur_o    : out    vl_logic;
        err_tlp_ur_lock_o: out    vl_logic;
        err_tlp_uc_o    : out    vl_logic;
        err_tlp_malformed_o: out    vl_logic;
        stat_tlp_cpl_ep_o: out    vl_logic;
        stat_tlp_cpl_abort_o: out    vl_logic;
        stat_tlp_cpl_ur_o: out    vl_logic;
        stat_tlp_ep_o   : out    vl_logic;
        check_raddr_o   : out    vl_logic_vector(63 downto 0);
        check_mem32_o   : out    vl_logic;
        check_mem64_o   : out    vl_logic;
        check_rio_o     : out    vl_logic;
        check_rdev_o    : out    vl_logic;
        check_rbus_o    : out    vl_logic;
        check_rfun_o    : out    vl_logic;
        check_rhit_i    : in     vl_logic;
        check_rhit_bar_i: in     vl_logic_vector;
        max_payload_i   : in     vl_logic_vector(2 downto 0);
        rhit_bar_lat3_i : in     vl_logic;
        legacy_mode_i   : in     vl_logic;
        legacy_cfg_access_i: in     vl_logic;
        ext_cfg_access_i: in     vl_logic;
        hotplug_msg_enable_i: in     vl_logic;
        td_ecrc_trim_i  : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DW : constant is 1;
    attribute mti_svvh_generic_type of FCW : constant is 1;
    attribute mti_svvh_generic_type of BARW : constant is 1;
    attribute mti_svvh_generic_type of DOWNSTREAM_PORT : constant is 1;
    attribute mti_svvh_generic_type of MPS : constant is 1;
    attribute mti_svvh_generic_type of TYPE1_UR : constant is 1;
end tlm_rx_data_snk;
