library verilog;
use verilog.vl_types.all;
entity mmureg_sv_unit is
end mmureg_sv_unit;
