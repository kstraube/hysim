library verilog;
use verilog.vl_types.all;
entity mmuwalk_sv_unit is
end mmuwalk_sv_unit;
