library verilog;
use verilog.vl_types.all;
entity libdebug is
end libdebug;
