library verilog;
use verilog.vl_types.all;
entity mac_gmii_sv_unit is
end mac_gmii_sv_unit;
