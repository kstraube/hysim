library verilog;
use verilog.vl_types.all;
entity libstd is
end libstd;
