library verilog;
use verilog.vl_types.all;
entity ddr2memctrl_fast_sv_unit is
end ddr2memctrl_fast_sv_unit;
