library verilog;
use verilog.vl_types.all;
entity libtm_cache_sv_unit is
end libtm_cache_sv_unit;
