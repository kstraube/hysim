library verilog;
use verilog.vl_types.all;
entity libopcodes is
end libopcodes;
