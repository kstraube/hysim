library verilog;
use verilog.vl_types.all;
entity pcie_blk_ll_credit is
    generic(
        C_STREAMING     : integer := 0;
        C_CALENDAR_STREAMING: integer := 4;
        C_CALENDAR_LEN  : integer := 9;
        C_CALENDAR_SUB_LEN: integer := 12;
        C_CALENDAR_SEQ  : vl_logic_vector(0 to 71) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        C_CALENDAR_SUB_SEQ: vl_logic_vector(0 to 95) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        MPS             : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        LEGACY_EP       : integer := 0;
        BFM_INIT_FC_PH  : integer := 0;
        BFM_INIT_FC_PD  : integer := 0;
        BFM_INIT_FC_NPH : integer := 0;
        BFM_INIT_FC_NPD : integer := 0;
        BFM_INIT_FC_CPLH: integer := 0;
        BFM_INIT_FC_CPLD: integer := 0
    );
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        mgmt_stats_credit_sel: out    vl_logic_vector(6 downto 0);
        mgmt_stats_credit: in     vl_logic_vector(11 downto 0);
        trn_pfc_ph_cl   : out    vl_logic_vector(7 downto 0);
        trn_pfc_nph_cl  : out    vl_logic_vector(7 downto 0);
        trn_pfc_cplh_cl : out    vl_logic_vector(7 downto 0);
        trn_pfc_cplh_cl_upd: out    vl_logic;
        trn_pfc_pd_cl   : out    vl_logic_vector(11 downto 0);
        trn_pfc_npd_cl  : out    vl_logic_vector(11 downto 0);
        trn_pfc_cpld_cl : out    vl_logic_vector(11 downto 0);
        trn_lnk_up_n    : in     vl_logic;
        trn_rfc_ph_av   : out    vl_logic_vector(7 downto 0);
        trn_rfc_pd_av   : out    vl_logic_vector(11 downto 0);
        trn_rfc_nph_av  : out    vl_logic_vector(7 downto 0);
        trn_rfc_npd_av  : out    vl_logic_vector(11 downto 0);
        trn_rfc_cplh_av : out    vl_logic_vector(7 downto 0);
        trn_rfc_cpld_av : out    vl_logic_vector(11 downto 0);
        trn_rcpl_streaming_n: in     vl_logic;
        rx_ch_credits_received: out    vl_logic_vector(7 downto 0);
        rx_ch_credits_received_inc: out    vl_logic;
        tx_ch_credits_consumed: out    vl_logic_vector(7 downto 0);
        tx_pd_credits_available: out    vl_logic_vector(11 downto 0);
        tx_pd_credits_consumed: out    vl_logic_vector(11 downto 0);
        tx_npd_credits_available: out    vl_logic_vector(11 downto 0);
        tx_npd_credits_consumed: out    vl_logic_vector(11 downto 0);
        tx_cd_credits_available: out    vl_logic_vector(11 downto 0);
        tx_cd_credits_consumed: out    vl_logic_vector(11 downto 0);
        clear_cpl_count : in     vl_logic;
        pd_credit_limited: out    vl_logic;
        npd_credit_limited: out    vl_logic;
        cd_credit_limited: out    vl_logic;
        l0_stats_cfg_transmitted: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of C_STREAMING : constant is 1;
    attribute mti_svvh_generic_type of C_CALENDAR_STREAMING : constant is 1;
    attribute mti_svvh_generic_type of C_CALENDAR_LEN : constant is 1;
    attribute mti_svvh_generic_type of C_CALENDAR_SUB_LEN : constant is 1;
    attribute mti_svvh_generic_type of C_CALENDAR_SEQ : constant is 1;
    attribute mti_svvh_generic_type of C_CALENDAR_SUB_SEQ : constant is 1;
    attribute mti_svvh_generic_type of MPS : constant is 1;
    attribute mti_svvh_generic_type of LEGACY_EP : constant is 1;
    attribute mti_svvh_generic_type of BFM_INIT_FC_PH : constant is 1;
    attribute mti_svvh_generic_type of BFM_INIT_FC_PD : constant is 1;
    attribute mti_svvh_generic_type of BFM_INIT_FC_NPH : constant is 1;
    attribute mti_svvh_generic_type of BFM_INIT_FC_NPD : constant is 1;
    attribute mti_svvh_generic_type of BFM_INIT_FC_CPLH : constant is 1;
    attribute mti_svvh_generic_type of BFM_INIT_FC_CPLD : constant is 1;
end pcie_blk_ll_credit;
