library verilog;
use verilog.vl_types.all;
entity dmmu_sv_unit is
end dmmu_sv_unit;
