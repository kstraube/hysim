library verilog;
use verilog.vl_types.all;
entity sim_memctrl_sv_unit is
end sim_memctrl_sv_unit;
