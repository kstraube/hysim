library verilog;
use verilog.vl_types.all;
entity techmap_sv_unit is
end techmap_sv_unit;
