library verilog;
use verilog.vl_types.all;
entity libmmu is
end libmmu;
