library verilog;
use verilog.vl_types.all;
entity tm_cpu_1ipc_sv_unit is
end tm_cpu_1ipc_sv_unit;
