library verilog;
use verilog.vl_types.all;
entity eth_cpu_control_sv_unit is
end eth_cpu_control_sv_unit;
