library verilog;
use verilog.vl_types.all;
entity dcacheram_sv_unit is
end dcacheram_sv_unit;
