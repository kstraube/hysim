library verilog;
use verilog.vl_types.all;
entity libtm_cache is
end libtm_cache;
