library verilog;
use verilog.vl_types.all;
entity memory_mmu_sv_unit is
end memory_mmu_sv_unit;
