library verilog;
use verilog.vl_types.all;
entity libmemif is
end libmemif;
