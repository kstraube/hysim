library verilog;
use verilog.vl_types.all;
entity dmabuf_sv_unit is
end dmabuf_sv_unit;
