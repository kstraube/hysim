library verilog;
use verilog.vl_types.all;
entity dramctrl_bee3_sv_unit is
end dramctrl_bee3_sv_unit;
