library verilog;
use verilog.vl_types.all;
entity disasm_sv_unit is
end disasm_sv_unit;
