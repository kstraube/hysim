library verilog;
use verilog.vl_types.all;
entity libeth is
end libeth;
