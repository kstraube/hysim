library verilog;
use verilog.vl_types.all;
entity clkrst_gen_sv_unit is
end clkrst_gen_sv_unit;
