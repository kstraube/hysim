library verilog;
use verilog.vl_types.all;
entity eth_dma_controller_sv_unit is
end eth_dma_controller_sv_unit;
