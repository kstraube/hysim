library verilog;
use verilog.vl_types.all;
entity dram_clkgen_sv_unit is
end dram_clkgen_sv_unit;
