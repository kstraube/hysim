library verilog;
use verilog.vl_types.all;
entity pcie_ep_top is
    generic(
        G_USER_RESETS   : integer := 0;
        G_SIM           : integer := 0;
        G_CHIPSCOPE     : integer := 0;
        INTF_CLK_FREQ   : integer := 0;
        REF_CLK_FREQ    : integer := 1;
        USE_V5FXT       : integer := 0;
        VEN_ID          : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0);
        DEV_ID          : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        REV_ID          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLASS_CODE      : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR0            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        BAR1            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR2            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        BAR3            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        BAR4            : integer := 0;
        BAR5            : integer := 0;
        CARDBUS_CIS_PTR : integer := 0;
        SUBSYS_VEN_ID   : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0);
        SUBSYS_ID       : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        XROM_BAR        : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        INTR_MSG_NUM    : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        SLT_IMPL        : vl_logic := Hi0;
        DEV_PORT_TYPE   : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        CAP_VER         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        CAPT_SLT_PWR_LIM_SC: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        CAPT_SLT_PWR_LIM_VA: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PWR_INDI_PRSNT  : vl_logic := Hi0;
        ATTN_INDI_PRSNT : vl_logic := Hi0;
        ATTN_BUTN_PRSNT : vl_logic := Hi0;
        EP_L1_ACCPT_LAT : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        EP_L0s_ACCPT_LAT: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        EXT_TAG_FLD_SUP : vl_logic := Hi0;
        PHANTM_FUNC_SUP : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        MPS             : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        L1_EXIT_LAT     : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        L0s_EXIT_LAT    : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        ASPM_SUP        : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        MAX_LNK_WDT     : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        MAX_LNK_SPD     : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        TRM_TLP_DGST_ECRC: vl_logic := Hi0;
        FRCE_NOSCRMBL   : vl_logic := Hi0;
        INFINITECOMPLETIONS: string  := "TRUE";
        VC0_CREDITS_PH  : integer := 8;
        VC0_CREDITS_NPH : integer := 8;
        CPL_STREAMING_PRIORITIZE_P_NP: integer := 0;
        SLOT_CLOCK_CONFIG: string  := "FALSE";
        C_CALENDAR_LEN  : vl_notype;
        C_CALENDAR_SEQ  : vl_notype;
        C_CALENDAR_SUB_LEN: integer := 12;
        C_CALENDAR_SUB_SEQ: vl_logic_vector(0 to 95) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        TX_DATACREDIT_FIX_EN: integer := 1;
        TX_DATACREDIT_FIX_1DWONLY: integer := 1;
        TX_DATACREDIT_FIX_MARGIN: integer := 6;
        TX_CPL_STALL_THRESHOLD: integer := 6;
        PME_SUP         : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        D2_SUP          : vl_logic := Hi1;
        D1_SUP          : vl_logic := Hi1;
        AUX_CT          : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        DSI             : vl_logic := Hi0;
        PME_CLK         : vl_logic := Hi0;
        PM_CAP_VER      : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        MSI_VECTOR      : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        MSI_8BIT_EN     : vl_logic := Hi0;
        PWR_CON_D0_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        CON_SCL_FCTR_D0_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PWR_CON_D1_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        CON_SCL_FCTR_D1_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PWR_CON_D2_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        CON_SCL_FCTR_D2_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PWR_CON_D3_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        CON_SCL_FCTR_D3_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PWR_DIS_D0_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        DIS_SCL_FCTR_D0_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PWR_DIS_D1_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        DIS_SCL_FCTR_D1_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PWR_DIS_D2_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        DIS_SCL_FCTR_D2_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PWR_DIS_D3_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        DIS_SCL_FCTR_D3_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        TXDIFFBOOST     : string  := "FALSE";
        GTDEBUGPORTS    : integer := 0
    );
    port(
        sys_clk         : in     vl_logic;
        sys_reset_n     : in     vl_logic;
        pci_exp_rxn     : in     vl_logic_vector;
        pci_exp_rxp     : in     vl_logic_vector;
        pci_exp_txn     : out    vl_logic_vector;
        pci_exp_txp     : out    vl_logic_vector;
        cfg_do          : out    vl_logic_vector(31 downto 0);
        cfg_di          : in     vl_logic_vector(31 downto 0);
        cfg_byte_en_n   : in     vl_logic_vector(3 downto 0);
        cfg_dwaddr      : in     vl_logic_vector(9 downto 0);
        cfg_rd_wr_done_n: out    vl_logic;
        cfg_wr_en_n     : in     vl_logic;
        cfg_rd_en_n     : in     vl_logic;
        cfg_err_cor_n   : in     vl_logic;
        cfg_err_ur_n    : in     vl_logic;
        cfg_err_ecrc_n  : in     vl_logic;
        cfg_err_cpl_timeout_n: in     vl_logic;
        cfg_err_cpl_abort_n: in     vl_logic;
        cfg_err_cpl_unexpect_n: in     vl_logic;
        cfg_err_posted_n: in     vl_logic;
        cfg_err_locked_n: in     vl_logic;
        cfg_interrupt_n : in     vl_logic;
        cfg_interrupt_rdy_n: out    vl_logic;
        cfg_interrupt_assert_n: in     vl_logic;
        cfg_interrupt_di: in     vl_logic_vector(7 downto 0);
        cfg_interrupt_do: out    vl_logic_vector(7 downto 0);
        cfg_interrupt_mmenable: out    vl_logic_vector(2 downto 0);
        cfg_interrupt_msienable: out    vl_logic;
        cfg_turnoff_ok_n: in     vl_logic;
        cfg_to_turnoff_n: out    vl_logic;
        cfg_pm_wake_n   : in     vl_logic;
        cfg_err_tlp_cpl_header: in     vl_logic_vector(47 downto 0);
        cfg_err_cpl_rdy_n: out    vl_logic;
        cfg_dsn         : in     vl_logic_vector(63 downto 0);
        cfg_trn_pending_n: in     vl_logic;
        cfg_status      : out    vl_logic_vector(15 downto 0);
        cfg_command     : out    vl_logic_vector(15 downto 0);
        cfg_dstatus     : out    vl_logic_vector(15 downto 0);
        cfg_dcommand    : out    vl_logic_vector(15 downto 0);
        cfg_lstatus     : out    vl_logic_vector(15 downto 0);
        cfg_lcommand    : out    vl_logic_vector(15 downto 0);
        cfg_bus_number  : out    vl_logic_vector(7 downto 0);
        cfg_device_number: out    vl_logic_vector(4 downto 0);
        cfg_function_number: out    vl_logic_vector(2 downto 0);
        cfg_pcie_link_state_n: out    vl_logic_vector(2 downto 0);
        trn_td          : in     vl_logic_vector(63 downto 0);
        trn_trem_n      : in     vl_logic_vector(7 downto 0);
        trn_tsof_n      : in     vl_logic;
        trn_teof_n      : in     vl_logic;
        trn_tsrc_rdy_n  : in     vl_logic;
        trn_tsrc_dsc_n  : in     vl_logic;
        trn_terrfwd_n   : in     vl_logic;
        trn_tdst_rdy_n  : out    vl_logic;
        trn_tdst_dsc_n  : out    vl_logic;
        trn_tbuf_av     : out    vl_logic_vector(3 downto 0);
        trn_rnp_ok_n    : in     vl_logic;
        trn_rdst_rdy_n  : in     vl_logic;
        trn_rd          : out    vl_logic_vector(63 downto 0);
        trn_rrem_n      : out    vl_logic_vector(7 downto 0);
        trn_rsof_n      : out    vl_logic;
        trn_reof_n      : out    vl_logic;
        trn_rsrc_rdy_n  : out    vl_logic;
        trn_rsrc_dsc_n  : out    vl_logic;
        trn_rerrfwd_n   : out    vl_logic;
        trn_rbar_hit_n  : out    vl_logic_vector(6 downto 0);
        trn_rfc_nph_av  : out    vl_logic_vector(7 downto 0);
        trn_rfc_npd_av  : out    vl_logic_vector(11 downto 0);
        trn_rfc_ph_av   : out    vl_logic_vector(7 downto 0);
        trn_rfc_pd_av   : out    vl_logic_vector(11 downto 0);
        trn_rfc_cplh_av : out    vl_logic_vector(7 downto 0);
        trn_rfc_cpld_av : out    vl_logic_vector(11 downto 0);
        trn_rcpl_streaming_n: in     vl_logic;
        refclkout       : out    vl_logic;
        gt_dclk         : in     vl_logic;
        gt_daddr        : in     vl_logic_vector;
        gt_den          : in     vl_logic_vector;
        gt_dwen         : in     vl_logic_vector;
        gt_di           : in     vl_logic_vector;
        gt_do           : out    vl_logic_vector;
        gt_drdy         : out    vl_logic_vector;
        gt_txdiffctrl_0 : in     vl_logic_vector(2 downto 0);
        gt_txdiffctrl_1 : in     vl_logic_vector(2 downto 0);
        gt_txbuffctrl_0 : in     vl_logic_vector(2 downto 0);
        gt_txbuffctrl_1 : in     vl_logic_vector(2 downto 0);
        gt_txpreemphesis_0: in     vl_logic_vector(2 downto 0);
        gt_txpreemphesis_1: in     vl_logic_vector(2 downto 0);
        trn_clk         : out    vl_logic;
        trn_reset_n     : out    vl_logic;
        trn_lnk_up_n    : out    vl_logic;
        fast_train_simulation_only: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of G_USER_RESETS : constant is 1;
    attribute mti_svvh_generic_type of G_SIM : constant is 1;
    attribute mti_svvh_generic_type of G_CHIPSCOPE : constant is 1;
    attribute mti_svvh_generic_type of INTF_CLK_FREQ : constant is 1;
    attribute mti_svvh_generic_type of REF_CLK_FREQ : constant is 1;
    attribute mti_svvh_generic_type of USE_V5FXT : constant is 1;
    attribute mti_svvh_generic_type of VEN_ID : constant is 1;
    attribute mti_svvh_generic_type of DEV_ID : constant is 1;
    attribute mti_svvh_generic_type of REV_ID : constant is 1;
    attribute mti_svvh_generic_type of CLASS_CODE : constant is 1;
    attribute mti_svvh_generic_type of BAR0 : constant is 1;
    attribute mti_svvh_generic_type of BAR1 : constant is 1;
    attribute mti_svvh_generic_type of BAR2 : constant is 1;
    attribute mti_svvh_generic_type of BAR3 : constant is 1;
    attribute mti_svvh_generic_type of BAR4 : constant is 1;
    attribute mti_svvh_generic_type of BAR5 : constant is 1;
    attribute mti_svvh_generic_type of CARDBUS_CIS_PTR : constant is 1;
    attribute mti_svvh_generic_type of SUBSYS_VEN_ID : constant is 1;
    attribute mti_svvh_generic_type of SUBSYS_ID : constant is 1;
    attribute mti_svvh_generic_type of XROM_BAR : constant is 1;
    attribute mti_svvh_generic_type of INTR_MSG_NUM : constant is 1;
    attribute mti_svvh_generic_type of SLT_IMPL : constant is 1;
    attribute mti_svvh_generic_type of DEV_PORT_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CAP_VER : constant is 1;
    attribute mti_svvh_generic_type of CAPT_SLT_PWR_LIM_SC : constant is 1;
    attribute mti_svvh_generic_type of CAPT_SLT_PWR_LIM_VA : constant is 1;
    attribute mti_svvh_generic_type of PWR_INDI_PRSNT : constant is 1;
    attribute mti_svvh_generic_type of ATTN_INDI_PRSNT : constant is 1;
    attribute mti_svvh_generic_type of ATTN_BUTN_PRSNT : constant is 1;
    attribute mti_svvh_generic_type of EP_L1_ACCPT_LAT : constant is 1;
    attribute mti_svvh_generic_type of EP_L0s_ACCPT_LAT : constant is 1;
    attribute mti_svvh_generic_type of EXT_TAG_FLD_SUP : constant is 1;
    attribute mti_svvh_generic_type of PHANTM_FUNC_SUP : constant is 1;
    attribute mti_svvh_generic_type of MPS : constant is 1;
    attribute mti_svvh_generic_type of L1_EXIT_LAT : constant is 1;
    attribute mti_svvh_generic_type of L0s_EXIT_LAT : constant is 1;
    attribute mti_svvh_generic_type of ASPM_SUP : constant is 1;
    attribute mti_svvh_generic_type of MAX_LNK_WDT : constant is 1;
    attribute mti_svvh_generic_type of MAX_LNK_SPD : constant is 1;
    attribute mti_svvh_generic_type of TRM_TLP_DGST_ECRC : constant is 1;
    attribute mti_svvh_generic_type of FRCE_NOSCRMBL : constant is 1;
    attribute mti_svvh_generic_type of INFINITECOMPLETIONS : constant is 1;
    attribute mti_svvh_generic_type of VC0_CREDITS_PH : constant is 1;
    attribute mti_svvh_generic_type of VC0_CREDITS_NPH : constant is 1;
    attribute mti_svvh_generic_type of CPL_STREAMING_PRIORITIZE_P_NP : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CLOCK_CONFIG : constant is 1;
    attribute mti_svvh_generic_type of C_CALENDAR_LEN : constant is 3;
    attribute mti_svvh_generic_type of C_CALENDAR_SEQ : constant is 3;
    attribute mti_svvh_generic_type of C_CALENDAR_SUB_LEN : constant is 1;
    attribute mti_svvh_generic_type of C_CALENDAR_SUB_SEQ : constant is 1;
    attribute mti_svvh_generic_type of TX_DATACREDIT_FIX_EN : constant is 1;
    attribute mti_svvh_generic_type of TX_DATACREDIT_FIX_1DWONLY : constant is 1;
    attribute mti_svvh_generic_type of TX_DATACREDIT_FIX_MARGIN : constant is 1;
    attribute mti_svvh_generic_type of TX_CPL_STALL_THRESHOLD : constant is 1;
    attribute mti_svvh_generic_type of PME_SUP : constant is 1;
    attribute mti_svvh_generic_type of D2_SUP : constant is 1;
    attribute mti_svvh_generic_type of D1_SUP : constant is 1;
    attribute mti_svvh_generic_type of AUX_CT : constant is 1;
    attribute mti_svvh_generic_type of DSI : constant is 1;
    attribute mti_svvh_generic_type of PME_CLK : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_VER : constant is 1;
    attribute mti_svvh_generic_type of MSI_VECTOR : constant is 1;
    attribute mti_svvh_generic_type of MSI_8BIT_EN : constant is 1;
    attribute mti_svvh_generic_type of PWR_CON_D0_STATE : constant is 1;
    attribute mti_svvh_generic_type of CON_SCL_FCTR_D0_STATE : constant is 1;
    attribute mti_svvh_generic_type of PWR_CON_D1_STATE : constant is 1;
    attribute mti_svvh_generic_type of CON_SCL_FCTR_D1_STATE : constant is 1;
    attribute mti_svvh_generic_type of PWR_CON_D2_STATE : constant is 1;
    attribute mti_svvh_generic_type of CON_SCL_FCTR_D2_STATE : constant is 1;
    attribute mti_svvh_generic_type of PWR_CON_D3_STATE : constant is 1;
    attribute mti_svvh_generic_type of CON_SCL_FCTR_D3_STATE : constant is 1;
    attribute mti_svvh_generic_type of PWR_DIS_D0_STATE : constant is 1;
    attribute mti_svvh_generic_type of DIS_SCL_FCTR_D0_STATE : constant is 1;
    attribute mti_svvh_generic_type of PWR_DIS_D1_STATE : constant is 1;
    attribute mti_svvh_generic_type of DIS_SCL_FCTR_D1_STATE : constant is 1;
    attribute mti_svvh_generic_type of PWR_DIS_D2_STATE : constant is 1;
    attribute mti_svvh_generic_type of DIS_SCL_FCTR_D2_STATE : constant is 1;
    attribute mti_svvh_generic_type of PWR_DIS_D3_STATE : constant is 1;
    attribute mti_svvh_generic_type of DIS_SCL_FCTR_D3_STATE : constant is 1;
    attribute mti_svvh_generic_type of TXDIFFBOOST : constant is 1;
    attribute mti_svvh_generic_type of GTDEBUGPORTS : constant is 1;
end pcie_ep_top;
