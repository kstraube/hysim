library verilog;
use verilog.vl_types.all;
entity pcie_blk_plus_ll_rx is
    generic(
        BAR0            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        BAR1            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR2            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        BAR3            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        BAR4            : integer := 0;
        BAR5            : integer := 0;
        XROM_BAR        : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        MPS             : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        LEGACY_EP       : vl_logic := Hi0;
        TRIM_ECRC       : vl_logic := Hi0;
        CPL_STREAMING_PRIORITIZE_P_NP: integer := 0
    );
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        llk_rx_dst_req_n: out    vl_logic;
        llk_rx_dst_cont_req_n: out    vl_logic;
        llk_rx_ch_tc    : out    vl_logic_vector(2 downto 0);
        llk_rx_ch_fifo  : out    vl_logic_vector(1 downto 0);
        llk_tc_status   : in     vl_logic_vector(7 downto 0);
        llk_rx_data     : in     vl_logic_vector(63 downto 0);
        llk_rx_data_d   : out    vl_logic_vector(63 downto 0);
        llk_rx_src_rdy_n: in     vl_logic;
        llk_rx_src_last_req_n: in     vl_logic;
        llk_rx_src_dsc_n: in     vl_logic;
        llk_rx_sof_n    : in     vl_logic;
        llk_rx_eof_n    : in     vl_logic;
        llk_rx_valid_n  : in     vl_logic_vector(1 downto 0);
        llk_rx_ch_posted_available_n: in     vl_logic_vector(7 downto 0);
        llk_rx_ch_non_posted_available_n: in     vl_logic_vector(7 downto 0);
        llk_rx_ch_completion_available_n: in     vl_logic_vector(7 downto 0);
        llk_rx_preferred_type: in     vl_logic_vector(15 downto 0);
        trn_rd          : out    vl_logic_vector(63 downto 0);
        trn_rrem_n      : out    vl_logic_vector(7 downto 0);
        trn_rsof_n      : out    vl_logic;
        trn_reof_n      : out    vl_logic;
        trn_rsrc_rdy_n  : out    vl_logic;
        trn_rsrc_dsc_n  : out    vl_logic;
        trn_rerrfwd_n   : out    vl_logic;
        trn_rbar_hit_n  : out    vl_logic_vector(6 downto 0);
        trn_lnk_up_n    : in     vl_logic;
        trn_rnp_ok_n    : in     vl_logic;
        trn_rdst_rdy_n  : in     vl_logic;
        trn_rcpl_streaming_n: in     vl_logic;
        cfg_rx_bar0     : in     vl_logic_vector(31 downto 0);
        cfg_rx_bar1     : in     vl_logic_vector(31 downto 0);
        cfg_rx_bar2     : in     vl_logic_vector(31 downto 0);
        cfg_rx_bar3     : in     vl_logic_vector(31 downto 0);
        cfg_rx_bar4     : in     vl_logic_vector(31 downto 0);
        cfg_rx_bar5     : in     vl_logic_vector(31 downto 0);
        cfg_rx_xrom     : in     vl_logic_vector(31 downto 0);
        cfg_bus_number  : in     vl_logic_vector(7 downto 0);
        cfg_device_number: in     vl_logic_vector(4 downto 0);
        cfg_function_number: in     vl_logic_vector(2 downto 0);
        cfg_dcommand    : in     vl_logic_vector(15 downto 0);
        cfg_pmcsr       : in     vl_logic_vector(15 downto 0);
        io_space_enable : in     vl_logic;
        mem_space_enable: in     vl_logic;
        max_payload_size: in     vl_logic_vector(2 downto 0);
        rx_err_cpl_abort_n: out    vl_logic;
        rx_err_cpl_ur_n : out    vl_logic;
        rx_err_cpl_ep_n : out    vl_logic;
        rx_err_ep_n     : out    vl_logic;
        err_tlp_cpl_header: out    vl_logic_vector(47 downto 0);
        err_tlp_p       : out    vl_logic;
        err_tlp_ur      : out    vl_logic;
        err_tlp_ur_lock : out    vl_logic;
        err_tlp_uc      : out    vl_logic;
        err_tlp_malformed: out    vl_logic;
        l0_stats_tlp_received: in     vl_logic;
        rx_ch_credits_received: in     vl_logic_vector(7 downto 0);
        rx_ch_credits_received_inc: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of BAR0 : constant is 1;
    attribute mti_svvh_generic_type of BAR1 : constant is 1;
    attribute mti_svvh_generic_type of BAR2 : constant is 1;
    attribute mti_svvh_generic_type of BAR3 : constant is 1;
    attribute mti_svvh_generic_type of BAR4 : constant is 1;
    attribute mti_svvh_generic_type of BAR5 : constant is 1;
    attribute mti_svvh_generic_type of XROM_BAR : constant is 1;
    attribute mti_svvh_generic_type of MPS : constant is 1;
    attribute mti_svvh_generic_type of LEGACY_EP : constant is 1;
    attribute mti_svvh_generic_type of TRIM_ECRC : constant is 1;
    attribute mti_svvh_generic_type of CPL_STREAMING_PRIORITIZE_P_NP : constant is 1;
end pcie_blk_plus_ll_rx;
