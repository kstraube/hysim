library verilog;
use verilog.vl_types.all;
entity memif_sv_unit is
end memif_sv_unit;
