library verilog;
use verilog.vl_types.all;
entity ddr2 is
    generic(
        TCK_MIN         : integer := 2500;
        TJIT_PER        : integer := 100;
        TJIT_DUTY       : integer := 100;
        TJIT_CC         : integer := 200;
        TERR_2PER       : integer := 150;
        TERR_3PER       : integer := 175;
        TERR_4PER       : integer := 200;
        TERR_5PER       : integer := 200;
        TERR_N1PER      : integer := 300;
        TERR_N2PER      : integer := 450;
        TQHS            : integer := 300;
        TAC             : integer := 400;
        TDS             : integer := 50;
        TDH             : integer := 125;
        TDQSCK          : integer := 350;
        TDQSQ           : integer := 200;
        TIS             : integer := 175;
        TIH             : integer := 250;
        TRC             : integer := 55000;
        TRCD            : integer := 15000;
        TWTR            : integer := 7500;
        TRP             : integer := 15000;
        TRPA            : integer := 17500;
        TXARDS          : integer := 8;
        TXARD           : integer := 2;
        TXP             : integer := 2;
        TANPD           : integer := 3;
        TAXPD           : integer := 10;
        CL_TIME         : integer := 15000;
        TFAW            : integer := 35000;
        AL_MIN          : integer := 0;
        AL_MAX          : integer := 6;
        CL_MIN          : integer := 3;
        CL_MAX          : integer := 7;
        WR_MIN          : integer := 2;
        WR_MAX          : integer := 8;
        BL_MIN          : integer := 4;
        BL_MAX          : integer := 8;
        TCK_MAX         : integer := 8000;
        TCH_MIN         : real    := 0.480000;
        TCH_MAX         : real    := 0.520000;
        TCL_MIN         : real    := 0.480000;
        TCL_MAX         : real    := 0.520000;
        TLZ             : vl_notype;
        THZ             : vl_notype;
        TDIPW           : real    := 0.350000;
        TDQSH           : real    := 0.350000;
        TDQSL           : real    := 0.350000;
        TDSS            : real    := 0.200000;
        TDSH            : real    := 0.200000;
        TWPRE           : real    := 0.350000;
        TWPST           : real    := 0.400000;
        TDQSS           : real    := 0.250000;
        TIPW            : real    := 0.600000;
        TCCD            : integer := 2;
        TRAS_MIN        : integer := 40000;
        TRAS_MAX        : integer := 70000000;
        TRTP            : integer := 7500;
        TWR             : integer := 15000;
        TMRD            : integer := 2;
        TDLLK           : integer := 200;
        TRFC_MIN        : integer := 127500;
        TRFC_MAX        : integer := 70000000;
        TXSNR           : vl_notype;
        TXSRD           : integer := 200;
        TISXR           : vl_notype;
        TAOND           : integer := 2;
        TAOFD           : real    := 2.500000;
        TAONPD          : integer := 2000;
        TAOFPD          : integer := 2000;
        TMOD            : integer := 12000;
        TCKE            : integer := 3;
        ADDR_BITS       : integer := 14;
        ROW_BITS        : integer := 14;
        COL_BITS        : integer := 10;
        DM_BITS         : integer := 1;
        DQ_BITS         : integer := 8;
        DQS_BITS        : integer := 1;
        TRRD            : integer := 7500;
        CS_BITS         : integer := 2;
        RANKS           : integer := 2;
        BA_BITS         : integer := 3;
        MEM_BITS        : integer := 22;
        AP              : integer := 10;
        BL_BITS         : integer := 3;
        BO_BITS         : integer := 2;
        STOP_ON_ERROR   : integer := 1;
        DEBUG           : integer := 0;
        BUS_DELAY       : integer := 6000;
        RANDOM_OUT_DELAY: integer := 0;
        RANDOM_SEED     : integer := 711689044;
        RDQSEN_PRE      : integer := 2;
        RDQSEN_PST      : integer := 1;
        RDQS_PRE        : integer := 2;
        RDQS_PST        : integer := 1;
        RDQEN_PRE       : integer := 0;
        RDQEN_PST       : integer := 0;
        WDQS_PRE        : integer := 1;
        WDQS_PST        : integer := 1;
        LOAD_MODE       : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        REFRESH         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        PRECHARGE       : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        ACTIVATE        : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        WRITE           : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        READ            : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        NOP             : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        PWR_DOWN        : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        SELF_REF        : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi1)
    );
    port(
        ck              : in     vl_logic;
        ck_n            : in     vl_logic;
        cke             : in     vl_logic;
        cs_n            : in     vl_logic;
        ras_n           : in     vl_logic;
        cas_n           : in     vl_logic;
        we_n            : in     vl_logic;
        dm_rdqs         : inout  vl_logic_vector;
        ba              : in     vl_logic_vector;
        addr            : in     vl_logic_vector;
        dq              : inout  vl_logic_vector;
        dqs             : inout  vl_logic_vector;
        dqs_n           : inout  vl_logic_vector;
        rdqs_n          : out    vl_logic_vector;
        odt             : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of TCK_MIN : constant is 1;
    attribute mti_svvh_generic_type of TJIT_PER : constant is 1;
    attribute mti_svvh_generic_type of TJIT_DUTY : constant is 1;
    attribute mti_svvh_generic_type of TJIT_CC : constant is 1;
    attribute mti_svvh_generic_type of TERR_2PER : constant is 1;
    attribute mti_svvh_generic_type of TERR_3PER : constant is 1;
    attribute mti_svvh_generic_type of TERR_4PER : constant is 1;
    attribute mti_svvh_generic_type of TERR_5PER : constant is 1;
    attribute mti_svvh_generic_type of TERR_N1PER : constant is 1;
    attribute mti_svvh_generic_type of TERR_N2PER : constant is 1;
    attribute mti_svvh_generic_type of TQHS : constant is 1;
    attribute mti_svvh_generic_type of TAC : constant is 1;
    attribute mti_svvh_generic_type of TDS : constant is 1;
    attribute mti_svvh_generic_type of TDH : constant is 1;
    attribute mti_svvh_generic_type of TDQSCK : constant is 1;
    attribute mti_svvh_generic_type of TDQSQ : constant is 1;
    attribute mti_svvh_generic_type of TIS : constant is 1;
    attribute mti_svvh_generic_type of TIH : constant is 1;
    attribute mti_svvh_generic_type of TRC : constant is 1;
    attribute mti_svvh_generic_type of TRCD : constant is 1;
    attribute mti_svvh_generic_type of TWTR : constant is 1;
    attribute mti_svvh_generic_type of TRP : constant is 1;
    attribute mti_svvh_generic_type of TRPA : constant is 1;
    attribute mti_svvh_generic_type of TXARDS : constant is 1;
    attribute mti_svvh_generic_type of TXARD : constant is 1;
    attribute mti_svvh_generic_type of TXP : constant is 1;
    attribute mti_svvh_generic_type of TANPD : constant is 1;
    attribute mti_svvh_generic_type of TAXPD : constant is 1;
    attribute mti_svvh_generic_type of CL_TIME : constant is 1;
    attribute mti_svvh_generic_type of TFAW : constant is 1;
    attribute mti_svvh_generic_type of AL_MIN : constant is 1;
    attribute mti_svvh_generic_type of AL_MAX : constant is 1;
    attribute mti_svvh_generic_type of CL_MIN : constant is 1;
    attribute mti_svvh_generic_type of CL_MAX : constant is 1;
    attribute mti_svvh_generic_type of WR_MIN : constant is 1;
    attribute mti_svvh_generic_type of WR_MAX : constant is 1;
    attribute mti_svvh_generic_type of BL_MIN : constant is 1;
    attribute mti_svvh_generic_type of BL_MAX : constant is 1;
    attribute mti_svvh_generic_type of TCK_MAX : constant is 1;
    attribute mti_svvh_generic_type of TCH_MIN : constant is 1;
    attribute mti_svvh_generic_type of TCH_MAX : constant is 1;
    attribute mti_svvh_generic_type of TCL_MIN : constant is 1;
    attribute mti_svvh_generic_type of TCL_MAX : constant is 1;
    attribute mti_svvh_generic_type of TLZ : constant is 3;
    attribute mti_svvh_generic_type of THZ : constant is 3;
    attribute mti_svvh_generic_type of TDIPW : constant is 1;
    attribute mti_svvh_generic_type of TDQSH : constant is 1;
    attribute mti_svvh_generic_type of TDQSL : constant is 1;
    attribute mti_svvh_generic_type of TDSS : constant is 1;
    attribute mti_svvh_generic_type of TDSH : constant is 1;
    attribute mti_svvh_generic_type of TWPRE : constant is 1;
    attribute mti_svvh_generic_type of TWPST : constant is 1;
    attribute mti_svvh_generic_type of TDQSS : constant is 1;
    attribute mti_svvh_generic_type of TIPW : constant is 1;
    attribute mti_svvh_generic_type of TCCD : constant is 1;
    attribute mti_svvh_generic_type of TRAS_MIN : constant is 1;
    attribute mti_svvh_generic_type of TRAS_MAX : constant is 1;
    attribute mti_svvh_generic_type of TRTP : constant is 1;
    attribute mti_svvh_generic_type of TWR : constant is 1;
    attribute mti_svvh_generic_type of TMRD : constant is 1;
    attribute mti_svvh_generic_type of TDLLK : constant is 1;
    attribute mti_svvh_generic_type of TRFC_MIN : constant is 1;
    attribute mti_svvh_generic_type of TRFC_MAX : constant is 1;
    attribute mti_svvh_generic_type of TXSNR : constant is 3;
    attribute mti_svvh_generic_type of TXSRD : constant is 1;
    attribute mti_svvh_generic_type of TISXR : constant is 3;
    attribute mti_svvh_generic_type of TAOND : constant is 1;
    attribute mti_svvh_generic_type of TAOFD : constant is 1;
    attribute mti_svvh_generic_type of TAONPD : constant is 1;
    attribute mti_svvh_generic_type of TAOFPD : constant is 1;
    attribute mti_svvh_generic_type of TMOD : constant is 1;
    attribute mti_svvh_generic_type of TCKE : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BITS : constant is 1;
    attribute mti_svvh_generic_type of ROW_BITS : constant is 1;
    attribute mti_svvh_generic_type of COL_BITS : constant is 1;
    attribute mti_svvh_generic_type of DM_BITS : constant is 1;
    attribute mti_svvh_generic_type of DQ_BITS : constant is 1;
    attribute mti_svvh_generic_type of DQS_BITS : constant is 1;
    attribute mti_svvh_generic_type of TRRD : constant is 1;
    attribute mti_svvh_generic_type of CS_BITS : constant is 1;
    attribute mti_svvh_generic_type of RANKS : constant is 1;
    attribute mti_svvh_generic_type of BA_BITS : constant is 1;
    attribute mti_svvh_generic_type of MEM_BITS : constant is 1;
    attribute mti_svvh_generic_type of AP : constant is 1;
    attribute mti_svvh_generic_type of BL_BITS : constant is 1;
    attribute mti_svvh_generic_type of BO_BITS : constant is 1;
    attribute mti_svvh_generic_type of STOP_ON_ERROR : constant is 1;
    attribute mti_svvh_generic_type of DEBUG : constant is 1;
    attribute mti_svvh_generic_type of BUS_DELAY : constant is 1;
    attribute mti_svvh_generic_type of RANDOM_OUT_DELAY : constant is 1;
    attribute mti_svvh_generic_type of RANDOM_SEED : constant is 1;
    attribute mti_svvh_generic_type of RDQSEN_PRE : constant is 1;
    attribute mti_svvh_generic_type of RDQSEN_PST : constant is 1;
    attribute mti_svvh_generic_type of RDQS_PRE : constant is 1;
    attribute mti_svvh_generic_type of RDQS_PST : constant is 1;
    attribute mti_svvh_generic_type of RDQEN_PRE : constant is 1;
    attribute mti_svvh_generic_type of RDQEN_PST : constant is 1;
    attribute mti_svvh_generic_type of WDQS_PRE : constant is 1;
    attribute mti_svvh_generic_type of WDQS_PST : constant is 1;
    attribute mti_svvh_generic_type of LOAD_MODE : constant is 1;
    attribute mti_svvh_generic_type of REFRESH : constant is 1;
    attribute mti_svvh_generic_type of PRECHARGE : constant is 1;
    attribute mti_svvh_generic_type of ACTIVATE : constant is 1;
    attribute mti_svvh_generic_type of WRITE : constant is 1;
    attribute mti_svvh_generic_type of READ : constant is 1;
    attribute mti_svvh_generic_type of NOP : constant is 1;
    attribute mti_svvh_generic_type of PWR_DOWN : constant is 1;
    attribute mti_svvh_generic_type of SELF_REF : constant is 1;
end ddr2;
