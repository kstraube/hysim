library verilog;
use verilog.vl_types.all;
entity itlb_2way_split_sv_unit is
end itlb_2way_split_sv_unit;
