library verilog;
use verilog.vl_types.all;
entity icacheram_sv_unit is
end icacheram_sv_unit;
