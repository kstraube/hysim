library verilog;
use verilog.vl_types.all;
entity xalu_sv_unit is
end xalu_sv_unit;
