library verilog;
use verilog.vl_types.all;
entity aludiv_sv_unit is
end aludiv_sv_unit;
