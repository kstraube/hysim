library verilog;
use verilog.vl_types.all;
entity tm_cpu_none_sv_unit is
end tm_cpu_none_sv_unit;
