library verilog;
use verilog.vl_types.all;
entity libfp is
end libfp;
