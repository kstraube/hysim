library verilog;
use verilog.vl_types.all;
entity timer_sv_unit is
end timer_sv_unit;
