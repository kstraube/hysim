library verilog;
use verilog.vl_types.all;
entity sync_lutram_fifo_sv_unit is
end sync_lutram_fifo_sv_unit;
