library verilog;
use verilog.vl_types.all;
entity libiu is
end libiu;
