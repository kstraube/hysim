library verilog;
use verilog.vl_types.all;
entity pcie_top_wrapper is
    generic(
        G_SIM           : integer := 1;
        G_USER_RESETS   : integer := 0;
        REF_CLK_FREQ    : integer := 1;
        COMPONENTTYPE   : integer := 0;
        NO_OF_LANES     : integer := 1;
        CLKRATIO        : integer := 1;
        CLKDIVIDED      : string  := "FALSE";
        USE_V5FXT       : integer := 0;
        VENDORID        : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0);
        DEVICEID        : vl_logic_vector(0 to 15) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        REVISIONID      : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SUBSYSTEMVENDORID: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0);
        SUBSYSTEMID     : vl_logic_vector(0 to 15) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        CLASSCODE       : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CARDBUSCISPOINTER: integer := 0;
        INTERRUPTPIN    : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR0EXIST       : string  := "TRUE";
        BAR0IOMEMN      : integer := 0;
        BAR064          : integer := 0;
        BAR0PREFETCHABLE: string  := "FALSE";
        BAR0MASKWIDTH   : vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        BAR1EXIST       : string  := "FALSE";
        BAR1IOMEMN      : integer := 0;
        BAR1PREFETCHABLE: string  := "FALSE";
        BAR1MASKWIDTH   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR2EXIST       : string  := "FALSE";
        BAR2IOMEMN      : integer := 0;
        BAR264          : integer := 0;
        BAR2PREFETCHABLE: string  := "FALSE";
        BAR2MASKWIDTH   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR3EXIST       : string  := "FALSE";
        BAR3IOMEMN      : integer := 0;
        BAR3PREFETCHABLE: string  := "FALSE";
        BAR3MASKWIDTH   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR4EXIST       : string  := "FALSE";
        BAR4IOMEMN      : integer := 0;
        BAR464          : integer := 0;
        BAR4PREFETCHABLE: string  := "FALSE";
        BAR4MASKWIDTH   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR5EXIST       : string  := "FALSE";
        BAR5IOMEMN      : integer := 0;
        BAR5PREFETCHABLE: string  := "FALSE";
        BAR5MASKWIDTH   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        MAXPAYLOADSIZE  : integer := 0;
        DEVICECAPABILITYENDPOINTL0SLATENCY: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        DEVICECAPABILITYENDPOINTL1LATENCY: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        LINKCAPABILITYASPMSUPPORTEN: integer := 0;
        L0SEXITLATENCY  : integer := 7;
        L0SEXITLATENCYCOMCLK: integer := 7;
        L1EXITLATENCY   : integer := 7;
        L1EXITLATENCYCOMCLK: integer := 7;
        MSIENABLE       : integer := 0;
        DSNENABLE       : integer := 0;
        VCENABLE        : integer := 0;
        MSICAPABILITYMULTIMSGCAP: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PMCAPABILITYDSI : string  := "TRUE";
        PMCAPABILITYPMESUPPORT: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        PORTVCCAPABILITYEXTENDEDVCCOUNT: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PORTVCCAPABILITYVCARBCAP: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        LOWPRIORITYVCCOUNT: integer := 0;
        DEVICESERIALNUMBER: vl_logic_vector(0 to 63) := (Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1);
        FORCENOSCRAMBLING: vl_logic := Hi0;
        INFINITECOMPLETIONS: string  := "TRUE";
        VC0_CREDITS_PH  : integer := 8;
        VC0_CREDITS_NPH : integer := 8;
        LINKSTATUSSLOTCLOCKCONFIG: string  := "FALSE";
        TXTSNFTS        : integer := 255;
        TXTSNFTSCOMCLK  : integer := 255;
        RESETMODE       : string  := "TRUE";
        RETRYRAMSIZE    : integer := 9;
        VC0RXFIFOSIZEP  : integer := 1024;
        VC0RXFIFOSIZENP : integer := 192;
        VC0RXFIFOSIZEC  : integer := 1024;
        VC1RXFIFOSIZEP  : integer := 0;
        VC1RXFIFOSIZENP : integer := 0;
        VC1RXFIFOSIZEC  : integer := 0;
        VC0TXFIFOSIZEP  : integer := 1024;
        VC0TXFIFOSIZENP : integer := 192;
        VC0TXFIFOSIZEC  : integer := 1024;
        VC1TXFIFOSIZEP  : integer := 0;
        VC1TXFIFOSIZENP : integer := 0;
        VC1TXFIFOSIZEC  : integer := 0;
        TXDIFFBOOST     : string  := "FALSE";
        GTDEBUGPORTS    : integer := 0
    );
    port(
        user_reset_n    : in     vl_logic;
        core_clk        : out    vl_logic;
        user_clk        : out    vl_logic;
        clock_lock      : out    vl_logic;
        gsr             : in     vl_logic;
        crm_urst_n      : in     vl_logic;
        crm_nvrst_n     : in     vl_logic;
        crm_mgmt_rst_n  : in     vl_logic;
        crm_user_cfg_rst_n: in     vl_logic;
        crm_mac_rst_n   : in     vl_logic;
        crm_link_rst_n  : in     vl_logic;
        compliance_avoid: in     vl_logic;
        l0_cfg_loopback_master: in     vl_logic;
        l0_transactions_pending: in     vl_logic;
        l0_set_completer_abort_error: in     vl_logic;
        l0_set_detected_corr_error: in     vl_logic;
        l0_set_detected_fatal_error: in     vl_logic;
        l0_set_detected_nonfatal_error: in     vl_logic;
        l0_set_user_detected_parity_error: in     vl_logic;
        l0_set_user_master_data_parity: in     vl_logic;
        l0_set_user_received_master_abort: in     vl_logic;
        l0_set_user_received_target_abort: in     vl_logic;
        l0_set_user_system_error: in     vl_logic;
        l0_set_user_signalled_target_abort: in     vl_logic;
        l0_set_completion_timeout_uncorr_error: in     vl_logic;
        l0_set_completion_timeout_corr_error: in     vl_logic;
        l0_set_unexpected_completion_uncorr_error: in     vl_logic;
        l0_set_unexpected_completion_corr_error: in     vl_logic;
        l0_set_unsupported_request_nonposted_error: in     vl_logic;
        l0_set_unsupported_request_other_error: in     vl_logic;
        l0_legacy_int_funct0: in     vl_logic;
        l0_msi_request0 : in     vl_logic_vector(3 downto 0);
        mgmt_wdata      : in     vl_logic_vector(31 downto 0);
        mgmt_bwren      : in     vl_logic_vector(3 downto 0);
        mgmt_wren       : in     vl_logic;
        mgmt_addr       : in     vl_logic_vector(10 downto 0);
        mgmt_rden       : in     vl_logic;
        mgmt_stats_credit_sel: in     vl_logic_vector(6 downto 0);
        crm_do_hot_reset_n: out    vl_logic;
        crm_pwr_soft_reset_n: out    vl_logic;
        mgmt_rdata      : out    vl_logic_vector(31 downto 0);
        mgmt_pso        : out    vl_logic_vector(16 downto 0);
        mgmt_stats_credit: out    vl_logic_vector(11 downto 0);
        l0_first_cfg_write_occurred: out    vl_logic;
        l0_cfg_loopback_ack: out    vl_logic;
        l0_rx_mac_link_error: out    vl_logic_vector(1 downto 0);
        l0_mac_link_up  : out    vl_logic;
        l0_mac_negotiated_link_width: out    vl_logic_vector(3 downto 0);
        l0_mac_link_training: out    vl_logic;
        l0_ltssm_state  : out    vl_logic_vector(3 downto 0);
        l0_mac_new_state_ack: out    vl_logic;
        l0_mac_rx_l0s_state: out    vl_logic;
        l0_mac_entered_l0: out    vl_logic;
        l0_dl_up_down   : out    vl_logic_vector(7 downto 0);
        l0_dll_error_vector: out    vl_logic_vector(6 downto 0);
        l0_completer_id : out    vl_logic_vector(12 downto 0);
        l0_msi_enable0  : out    vl_logic;
        l0_multi_msg_en0: out    vl_logic_vector(2 downto 0);
        l0_stats_dllp_received: out    vl_logic;
        l0_stats_dllp_transmitted: out    vl_logic;
        l0_stats_os_received: out    vl_logic;
        l0_stats_os_transmitted: out    vl_logic;
        l0_stats_tlp_received: out    vl_logic;
        l0_stats_tlp_transmitted: out    vl_logic;
        l0_stats_cfg_received: out    vl_logic;
        l0_stats_cfg_transmitted: out    vl_logic;
        l0_stats_cfg_other_received: out    vl_logic;
        l0_stats_cfg_other_transmitted: out    vl_logic;
        l0_pwr_state0   : out    vl_logic_vector(1 downto 0);
        l0_pwr_l23_ready_state: out    vl_logic;
        l0_pwr_tx_l0s_state: out    vl_logic;
        l0_pwr_turn_off_req: out    vl_logic;
        l0_pme_req_in   : in     vl_logic;
        l0_pme_ack      : out    vl_logic;
        io_space_enable : out    vl_logic;
        mem_space_enable: out    vl_logic;
        bus_master_enable: out    vl_logic;
        parity_error_response: out    vl_logic;
        serr_enable     : out    vl_logic;
        interrupt_disable: out    vl_logic;
        ur_reporting_enable: out    vl_logic;
        llk_tx_data     : in     vl_logic_vector(63 downto 0);
        llk_tx_src_rdy_n: in     vl_logic;
        llk_tx_sof_n    : in     vl_logic;
        llk_tx_eof_n    : in     vl_logic;
        llk_tx_sop_n    : in     vl_logic;
        llk_tx_eop_n    : in     vl_logic;
        llk_tx_enable_n : in     vl_logic_vector(1 downto 0);
        llk_tx_ch_tc    : in     vl_logic_vector(2 downto 0);
        llk_tx_ch_fifo  : in     vl_logic_vector(1 downto 0);
        llk_tx_src_dsc_n: in     vl_logic;
        llk_tx_dst_rdy_n: out    vl_logic;
        llk_tx_chan_space: out    vl_logic_vector(9 downto 0);
        llk_tx_ch_posted_ready_n: out    vl_logic_vector(7 downto 0);
        llk_tx_ch_non_posted_ready_n: out    vl_logic_vector(7 downto 0);
        llk_tx_ch_completion_ready_n: out    vl_logic_vector(7 downto 0);
        llk_rx_dst_req_n: in     vl_logic;
        llk_rx_dst_cont_req_n: in     vl_logic;
        llk_rx_ch_tc    : in     vl_logic_vector(2 downto 0);
        llk_rx_ch_fifo  : in     vl_logic_vector(1 downto 0);
        llk_tc_status   : out    vl_logic_vector(7 downto 0);
        llk_rx_data     : out    vl_logic_vector(63 downto 0);
        llk_rx_src_rdy_n: out    vl_logic;
        llk_rx_src_last_req_n: out    vl_logic;
        llk_rx_sof_n    : out    vl_logic;
        llk_rx_eof_n    : out    vl_logic;
        llk_rx_sop_n    : out    vl_logic;
        llk_rx_eop_n    : out    vl_logic;
        llk_rx_valid_n  : out    vl_logic_vector(1 downto 0);
        llk_rx_ch_posted_available_n: out    vl_logic_vector(7 downto 0);
        llk_rx_ch_non_posted_available_n: out    vl_logic_vector(7 downto 0);
        llk_rx_ch_completion_available_n: out    vl_logic_vector(7 downto 0);
        llk_rx_preferred_type: out    vl_logic_vector(15 downto 0);
        RXN             : in     vl_logic_vector;
        RXP             : in     vl_logic_vector;
        TXN             : out    vl_logic_vector;
        TXP             : out    vl_logic_vector;
        GTPCLK_bufg     : out    vl_logic;
        REFCLKOUT_bufg  : out    vl_logic;
        PLLLKDET_OUT    : out    vl_logic_vector(3 downto 0);
        RESETDONE       : out    vl_logic_vector(7 downto 0);
        DEBUG           : out    vl_logic_vector(338 downto 0);
        GTPRESET        : in     vl_logic;
        REFCLK          : in     vl_logic;
        gt_rx_present   : in     vl_logic_vector(7 downto 0);
        gt_dclk         : in     vl_logic;
        gt_daddr        : in     vl_logic_vector;
        gt_den          : in     vl_logic_vector;
        gt_dwen         : in     vl_logic_vector;
        gt_di           : in     vl_logic_vector;
        gt_do           : out    vl_logic_vector;
        gt_drdy         : out    vl_logic_vector;
        gt_txdiffctrl_0 : in     vl_logic_vector(2 downto 0);
        gt_txdiffctrl_1 : in     vl_logic_vector(2 downto 0);
        gt_txbuffctrl_0 : in     vl_logic_vector(2 downto 0);
        gt_txbuffctrl_1 : in     vl_logic_vector(2 downto 0);
        gt_txpreemphesis_0: in     vl_logic_vector(2 downto 0);
        gt_txpreemphesis_1: in     vl_logic_vector(2 downto 0);
        trn_lnk_up_n    : in     vl_logic;
        max_payload_size: out    vl_logic_vector(2 downto 0);
        max_read_request_size: out    vl_logic_vector(2 downto 0);
        fast_train_simulation_only: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of G_SIM : constant is 1;
    attribute mti_svvh_generic_type of G_USER_RESETS : constant is 1;
    attribute mti_svvh_generic_type of REF_CLK_FREQ : constant is 1;
    attribute mti_svvh_generic_type of COMPONENTTYPE : constant is 1;
    attribute mti_svvh_generic_type of NO_OF_LANES : constant is 1;
    attribute mti_svvh_generic_type of CLKRATIO : constant is 1;
    attribute mti_svvh_generic_type of CLKDIVIDED : constant is 1;
    attribute mti_svvh_generic_type of USE_V5FXT : constant is 1;
    attribute mti_svvh_generic_type of VENDORID : constant is 1;
    attribute mti_svvh_generic_type of DEVICEID : constant is 1;
    attribute mti_svvh_generic_type of REVISIONID : constant is 1;
    attribute mti_svvh_generic_type of SUBSYSTEMVENDORID : constant is 1;
    attribute mti_svvh_generic_type of SUBSYSTEMID : constant is 1;
    attribute mti_svvh_generic_type of CLASSCODE : constant is 1;
    attribute mti_svvh_generic_type of CARDBUSCISPOINTER : constant is 1;
    attribute mti_svvh_generic_type of INTERRUPTPIN : constant is 2;
    attribute mti_svvh_generic_type of BAR0EXIST : constant is 1;
    attribute mti_svvh_generic_type of BAR0IOMEMN : constant is 1;
    attribute mti_svvh_generic_type of BAR064 : constant is 1;
    attribute mti_svvh_generic_type of BAR0PREFETCHABLE : constant is 1;
    attribute mti_svvh_generic_type of BAR0MASKWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR1EXIST : constant is 1;
    attribute mti_svvh_generic_type of BAR1IOMEMN : constant is 1;
    attribute mti_svvh_generic_type of BAR1PREFETCHABLE : constant is 1;
    attribute mti_svvh_generic_type of BAR1MASKWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR2EXIST : constant is 1;
    attribute mti_svvh_generic_type of BAR2IOMEMN : constant is 1;
    attribute mti_svvh_generic_type of BAR264 : constant is 1;
    attribute mti_svvh_generic_type of BAR2PREFETCHABLE : constant is 1;
    attribute mti_svvh_generic_type of BAR2MASKWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR3EXIST : constant is 1;
    attribute mti_svvh_generic_type of BAR3IOMEMN : constant is 1;
    attribute mti_svvh_generic_type of BAR3PREFETCHABLE : constant is 1;
    attribute mti_svvh_generic_type of BAR3MASKWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR4EXIST : constant is 1;
    attribute mti_svvh_generic_type of BAR4IOMEMN : constant is 1;
    attribute mti_svvh_generic_type of BAR464 : constant is 1;
    attribute mti_svvh_generic_type of BAR4PREFETCHABLE : constant is 1;
    attribute mti_svvh_generic_type of BAR4MASKWIDTH : constant is 2;
    attribute mti_svvh_generic_type of BAR5EXIST : constant is 1;
    attribute mti_svvh_generic_type of BAR5IOMEMN : constant is 1;
    attribute mti_svvh_generic_type of BAR5PREFETCHABLE : constant is 1;
    attribute mti_svvh_generic_type of BAR5MASKWIDTH : constant is 2;
    attribute mti_svvh_generic_type of MAXPAYLOADSIZE : constant is 1;
    attribute mti_svvh_generic_type of DEVICECAPABILITYENDPOINTL0SLATENCY : constant is 2;
    attribute mti_svvh_generic_type of DEVICECAPABILITYENDPOINTL1LATENCY : constant is 2;
    attribute mti_svvh_generic_type of LINKCAPABILITYASPMSUPPORTEN : constant is 1;
    attribute mti_svvh_generic_type of L0SEXITLATENCY : constant is 1;
    attribute mti_svvh_generic_type of L0SEXITLATENCYCOMCLK : constant is 1;
    attribute mti_svvh_generic_type of L1EXITLATENCY : constant is 1;
    attribute mti_svvh_generic_type of L1EXITLATENCYCOMCLK : constant is 1;
    attribute mti_svvh_generic_type of MSIENABLE : constant is 1;
    attribute mti_svvh_generic_type of DSNENABLE : constant is 1;
    attribute mti_svvh_generic_type of VCENABLE : constant is 1;
    attribute mti_svvh_generic_type of MSICAPABILITYMULTIMSGCAP : constant is 2;
    attribute mti_svvh_generic_type of PMCAPABILITYDSI : constant is 1;
    attribute mti_svvh_generic_type of PMCAPABILITYPMESUPPORT : constant is 1;
    attribute mti_svvh_generic_type of PORTVCCAPABILITYEXTENDEDVCCOUNT : constant is 2;
    attribute mti_svvh_generic_type of PORTVCCAPABILITYVCARBCAP : constant is 2;
    attribute mti_svvh_generic_type of LOWPRIORITYVCCOUNT : constant is 1;
    attribute mti_svvh_generic_type of DEVICESERIALNUMBER : constant is 1;
    attribute mti_svvh_generic_type of FORCENOSCRAMBLING : constant is 1;
    attribute mti_svvh_generic_type of INFINITECOMPLETIONS : constant is 1;
    attribute mti_svvh_generic_type of VC0_CREDITS_PH : constant is 1;
    attribute mti_svvh_generic_type of VC0_CREDITS_NPH : constant is 1;
    attribute mti_svvh_generic_type of LINKSTATUSSLOTCLOCKCONFIG : constant is 1;
    attribute mti_svvh_generic_type of TXTSNFTS : constant is 1;
    attribute mti_svvh_generic_type of TXTSNFTSCOMCLK : constant is 1;
    attribute mti_svvh_generic_type of RESETMODE : constant is 1;
    attribute mti_svvh_generic_type of RETRYRAMSIZE : constant is 1;
    attribute mti_svvh_generic_type of VC0RXFIFOSIZEP : constant is 1;
    attribute mti_svvh_generic_type of VC0RXFIFOSIZENP : constant is 1;
    attribute mti_svvh_generic_type of VC0RXFIFOSIZEC : constant is 1;
    attribute mti_svvh_generic_type of VC1RXFIFOSIZEP : constant is 1;
    attribute mti_svvh_generic_type of VC1RXFIFOSIZENP : constant is 1;
    attribute mti_svvh_generic_type of VC1RXFIFOSIZEC : constant is 1;
    attribute mti_svvh_generic_type of VC0TXFIFOSIZEP : constant is 1;
    attribute mti_svvh_generic_type of VC0TXFIFOSIZENP : constant is 1;
    attribute mti_svvh_generic_type of VC0TXFIFOSIZEC : constant is 1;
    attribute mti_svvh_generic_type of VC1TXFIFOSIZEP : constant is 1;
    attribute mti_svvh_generic_type of VC1TXFIFOSIZENP : constant is 1;
    attribute mti_svvh_generic_type of VC1TXFIFOSIZEC : constant is 1;
    attribute mti_svvh_generic_type of TXDIFFBOOST : constant is 1;
    attribute mti_svvh_generic_type of GTDEBUGPORTS : constant is 1;
end pcie_top_wrapper;
