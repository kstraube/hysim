library verilog;
use verilog.vl_types.all;
entity alumul_sv_unit is
end alumul_sv_unit;
