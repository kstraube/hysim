library verilog;
use verilog.vl_types.all;
entity dramif_sv_unit is
end dramif_sv_unit;
