library verilog;
use verilog.vl_types.all;
entity endpoint_blk_plus_v1_15 is
    generic(
        C_XDEVICE       : string  := "xc5vlx110t";
        USE_V5FXT       : integer := 0;
        PCI_EXP_LINK_WIDTH: integer := 1;
        PCI_EXP_INT_FREQ: integer := 0;
        PCI_EXP_REF_FREQ: integer := 0;
        PCI_EXP_TRN_DATA_WIDTH: integer := 64;
        PCI_EXP_TRN_REM_WIDTH: integer := 8;
        PCI_EXP_TRN_BUF_AV_WIDTH: integer := 4;
        PCI_EXP_BAR_HIT_WIDTH: integer := 7;
        PCI_EXP_FC_HDR_WIDTH: integer := 8;
        PCI_EXP_FC_DATA_WIDTH: integer := 12;
        PCI_EXP_CFG_DATA_WIDTH: integer := 32;
        PCI_EXP_CFG_ADDR_WIDTH: integer := 10;
        PCI_EXP_CFG_CPLHDR_WIDTH: integer := 48;
        PCI_EXP_CFG_BUSNUM_WIDTH: integer := 8;
        PCI_EXP_CFG_DEVNUM_WIDTH: integer := 5;
        PCI_EXP_CFG_FUNNUM_WIDTH: integer := 3;
        PCI_EXP_CFG_CAP_WIDTH: integer := 16;
        PCI_EXP_CFG_WIDTH: integer := 1024;
        VEN_ID_temp     : integer := 4334;
        VEN_ID          : vl_notype;
        DEV_ID          : vl_logic_vector(0 to 15) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        REV_ID          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLASS_CODE      : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR0            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR1            : integer := 0;
        BAR2            : integer := 0;
        BAR3            : integer := 0;
        BAR4            : integer := 0;
        BAR5            : integer := 0;
        CARDBUS_CIS_PTR : integer := 0;
        SUBSYS_VEN_ID_temp: integer := 4334;
        SUBSYS_ID_temp  : integer := 20560;
        SUBSYS_VEN_ID   : vl_notype;
        SUBSYS_ID       : vl_notype;
        XROM_BAR        : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        INTR_MSG_NUM    : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        SLT_IMPL        : integer := 0;
        DEV_PORT_TYPE   : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        CAP_VER         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        CAPT_SLT_PWR_LIM_SC: vl_logic_vector(0 to 1) := (Hi0, Hi0);
        CAPT_SLT_PWR_LIM_VA: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PWR_INDI_PRSNT  : integer := 0;
        ATTN_INDI_PRSNT : integer := 0;
        ATTN_BUTN_PRSNT : integer := 0;
        EP_L1_ACCPT_LAT : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        EP_L0s_ACCPT_LAT: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        EXT_TAG_FLD_SUP : integer := 1;
        PHANTM_FUNC_SUP : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        MPS             : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        L1_EXIT_LAT     : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        L0s_EXIT_LAT    : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        ASPM_SUP        : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        MAX_LNK_WDT     : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        MAX_LNK_SPD     : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        ACK_TO          : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        RPLY_TO         : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        MSI             : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        PCI_CONFIG_SPACE_ACCESS: integer := 0;
        EXT_CONFIG_SPACE_ACCESS: integer := 0;
        TRM_TLP_DGST_ECRC: integer := 0;
        FRCE_NOSCRMBL   : integer := 0;
        TWO_PLM_ATOCFGR : integer := 0;
        PME_SUP         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        D2_SUP          : integer := 0;
        D1_SUP          : integer := 0;
        AUX_CT          : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        DSI             : integer := 0;
        PME_CLK         : integer := 0;
        PM_CAP_VER      : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        PWR_CON_D0_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CON_SCL_FCTR_D0_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PWR_CON_D1_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CON_SCL_FCTR_D1_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PWR_CON_D2_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CON_SCL_FCTR_D2_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PWR_CON_D3_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CON_SCL_FCTR_D3_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PWR_DIS_D0_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DIS_SCL_FCTR_D0_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PWR_DIS_D1_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DIS_SCL_FCTR_D1_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PWR_DIS_D2_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DIS_SCL_FCTR_D2_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PWR_DIS_D3_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DIS_SCL_FCTR_D3_STATE: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CAL_BLK_DISABLE : integer := 0;
        SWAP_A_B_PAIRS  : integer := 0;
        INFINITECOMPLETIONS: string  := "TRUE";
        VC0_CREDITS_PH  : integer := 8;
        VC0_CREDITS_NPH : integer := 8;
        CPL_STREAMING_PRIORITIZE_P_NP: integer := 0;
        SLOT_CLK        : string  := "TRUE";
        TX_DIFF_BOOST   : string  := "TRUE";
        TXDIFFCTRL      : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        TXBUFDIFFCTRL   : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        TXPREEMPHASIS   : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        GT_Debug_Ports  : integer := 0;
        GTDEBUGPORTS    : integer := 0
    );
    port(
        pci_exp_txp     : out    vl_logic_vector;
        pci_exp_txn     : out    vl_logic_vector;
        pci_exp_rxp     : in     vl_logic_vector;
        pci_exp_rxn     : in     vl_logic_vector;
        trn_clk         : out    vl_logic;
        trn_reset_n     : out    vl_logic;
        trn_lnk_up_n    : out    vl_logic;
        trn_td          : in     vl_logic_vector;
        trn_trem_n      : in     vl_logic_vector;
        trn_tsof_n      : in     vl_logic;
        trn_teof_n      : in     vl_logic;
        trn_tsrc_rdy_n  : in     vl_logic;
        trn_tdst_rdy_n  : out    vl_logic;
        trn_tdst_dsc_n  : out    vl_logic;
        trn_tsrc_dsc_n  : in     vl_logic;
        trn_terrfwd_n   : in     vl_logic;
        trn_tbuf_av     : out    vl_logic_vector;
        trn_rd          : out    vl_logic_vector;
        trn_rrem_n      : out    vl_logic_vector;
        trn_rsof_n      : out    vl_logic;
        trn_reof_n      : out    vl_logic;
        trn_rsrc_rdy_n  : out    vl_logic;
        trn_rsrc_dsc_n  : out    vl_logic;
        trn_rdst_rdy_n  : in     vl_logic;
        trn_rerrfwd_n   : out    vl_logic;
        trn_rnp_ok_n    : in     vl_logic;
        trn_rbar_hit_n  : out    vl_logic_vector;
        trn_rfc_nph_av  : out    vl_logic_vector;
        trn_rfc_npd_av  : out    vl_logic_vector;
        trn_rfc_ph_av   : out    vl_logic_vector;
        trn_rfc_pd_av   : out    vl_logic_vector;
        trn_rcpl_streaming_n: in     vl_logic;
        cfg_do          : out    vl_logic_vector;
        cfg_rd_wr_done_n: out    vl_logic;
        cfg_di          : in     vl_logic_vector;
        cfg_byte_en_n   : in     vl_logic_vector;
        cfg_dwaddr      : in     vl_logic_vector;
        cfg_wr_en_n     : in     vl_logic;
        cfg_rd_en_n     : in     vl_logic;
        cfg_err_cor_n   : in     vl_logic;
        cfg_err_ur_n    : in     vl_logic;
        cfg_err_ecrc_n  : in     vl_logic;
        cfg_err_cpl_timeout_n: in     vl_logic;
        cfg_err_cpl_abort_n: in     vl_logic;
        cfg_err_cpl_unexpect_n: in     vl_logic;
        cfg_err_posted_n: in     vl_logic;
        cfg_err_tlp_cpl_header: in     vl_logic_vector;
        cfg_err_cpl_rdy_n: out    vl_logic;
        cfg_err_locked_n: in     vl_logic;
        cfg_interrupt_n : in     vl_logic;
        cfg_interrupt_rdy_n: out    vl_logic;
        cfg_interrupt_assert_n: in     vl_logic;
        cfg_interrupt_di: in     vl_logic_vector(7 downto 0);
        cfg_interrupt_do: out    vl_logic_vector(7 downto 0);
        cfg_interrupt_mmenable: out    vl_logic_vector(2 downto 0);
        cfg_interrupt_msienable: out    vl_logic;
        cfg_to_turnoff_n: out    vl_logic;
        cfg_pm_wake_n   : in     vl_logic;
        cfg_pcie_link_state_n: out    vl_logic_vector(2 downto 0);
        cfg_trn_pending_n: in     vl_logic;
        cfg_bus_number  : out    vl_logic_vector;
        cfg_device_number: out    vl_logic_vector;
        cfg_function_number: out    vl_logic_vector;
        cfg_dsn         : in     vl_logic_vector(63 downto 0);
        cfg_status      : out    vl_logic_vector;
        cfg_command     : out    vl_logic_vector;
        cfg_dstatus     : out    vl_logic_vector;
        cfg_dcommand    : out    vl_logic_vector;
        cfg_lstatus     : out    vl_logic_vector;
        cfg_lcommand    : out    vl_logic_vector;
        fast_train_simulation_only: in     vl_logic;
        sys_clk         : in     vl_logic;
        refclkout       : out    vl_logic;
        sys_reset_n     : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of C_XDEVICE : constant is 1;
    attribute mti_svvh_generic_type of USE_V5FXT : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_LINK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_INT_FREQ : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_REF_FREQ : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_TRN_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_TRN_REM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_TRN_BUF_AV_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_BAR_HIT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_FC_HDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_FC_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_CFG_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_CFG_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_CFG_CPLHDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_CFG_BUSNUM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_CFG_DEVNUM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_CFG_FUNNUM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_CFG_CAP_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXP_CFG_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of VEN_ID_temp : constant is 1;
    attribute mti_svvh_generic_type of VEN_ID : constant is 3;
    attribute mti_svvh_generic_type of DEV_ID : constant is 1;
    attribute mti_svvh_generic_type of REV_ID : constant is 1;
    attribute mti_svvh_generic_type of CLASS_CODE : constant is 1;
    attribute mti_svvh_generic_type of BAR0 : constant is 1;
    attribute mti_svvh_generic_type of BAR1 : constant is 1;
    attribute mti_svvh_generic_type of BAR2 : constant is 1;
    attribute mti_svvh_generic_type of BAR3 : constant is 1;
    attribute mti_svvh_generic_type of BAR4 : constant is 1;
    attribute mti_svvh_generic_type of BAR5 : constant is 1;
    attribute mti_svvh_generic_type of CARDBUS_CIS_PTR : constant is 1;
    attribute mti_svvh_generic_type of SUBSYS_VEN_ID_temp : constant is 1;
    attribute mti_svvh_generic_type of SUBSYS_ID_temp : constant is 1;
    attribute mti_svvh_generic_type of SUBSYS_VEN_ID : constant is 3;
    attribute mti_svvh_generic_type of SUBSYS_ID : constant is 3;
    attribute mti_svvh_generic_type of XROM_BAR : constant is 1;
    attribute mti_svvh_generic_type of INTR_MSG_NUM : constant is 1;
    attribute mti_svvh_generic_type of SLT_IMPL : constant is 1;
    attribute mti_svvh_generic_type of DEV_PORT_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CAP_VER : constant is 1;
    attribute mti_svvh_generic_type of CAPT_SLT_PWR_LIM_SC : constant is 1;
    attribute mti_svvh_generic_type of CAPT_SLT_PWR_LIM_VA : constant is 1;
    attribute mti_svvh_generic_type of PWR_INDI_PRSNT : constant is 1;
    attribute mti_svvh_generic_type of ATTN_INDI_PRSNT : constant is 1;
    attribute mti_svvh_generic_type of ATTN_BUTN_PRSNT : constant is 1;
    attribute mti_svvh_generic_type of EP_L1_ACCPT_LAT : constant is 1;
    attribute mti_svvh_generic_type of EP_L0s_ACCPT_LAT : constant is 1;
    attribute mti_svvh_generic_type of EXT_TAG_FLD_SUP : constant is 1;
    attribute mti_svvh_generic_type of PHANTM_FUNC_SUP : constant is 1;
    attribute mti_svvh_generic_type of MPS : constant is 1;
    attribute mti_svvh_generic_type of L1_EXIT_LAT : constant is 1;
    attribute mti_svvh_generic_type of L0s_EXIT_LAT : constant is 1;
    attribute mti_svvh_generic_type of ASPM_SUP : constant is 1;
    attribute mti_svvh_generic_type of MAX_LNK_WDT : constant is 1;
    attribute mti_svvh_generic_type of MAX_LNK_SPD : constant is 1;
    attribute mti_svvh_generic_type of ACK_TO : constant is 1;
    attribute mti_svvh_generic_type of RPLY_TO : constant is 1;
    attribute mti_svvh_generic_type of MSI : constant is 1;
    attribute mti_svvh_generic_type of PCI_CONFIG_SPACE_ACCESS : constant is 1;
    attribute mti_svvh_generic_type of EXT_CONFIG_SPACE_ACCESS : constant is 1;
    attribute mti_svvh_generic_type of TRM_TLP_DGST_ECRC : constant is 1;
    attribute mti_svvh_generic_type of FRCE_NOSCRMBL : constant is 1;
    attribute mti_svvh_generic_type of TWO_PLM_ATOCFGR : constant is 1;
    attribute mti_svvh_generic_type of PME_SUP : constant is 1;
    attribute mti_svvh_generic_type of D2_SUP : constant is 1;
    attribute mti_svvh_generic_type of D1_SUP : constant is 1;
    attribute mti_svvh_generic_type of AUX_CT : constant is 1;
    attribute mti_svvh_generic_type of DSI : constant is 1;
    attribute mti_svvh_generic_type of PME_CLK : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_VER : constant is 1;
    attribute mti_svvh_generic_type of PWR_CON_D0_STATE : constant is 1;
    attribute mti_svvh_generic_type of CON_SCL_FCTR_D0_STATE : constant is 1;
    attribute mti_svvh_generic_type of PWR_CON_D1_STATE : constant is 1;
    attribute mti_svvh_generic_type of CON_SCL_FCTR_D1_STATE : constant is 1;
    attribute mti_svvh_generic_type of PWR_CON_D2_STATE : constant is 1;
    attribute mti_svvh_generic_type of CON_SCL_FCTR_D2_STATE : constant is 1;
    attribute mti_svvh_generic_type of PWR_CON_D3_STATE : constant is 1;
    attribute mti_svvh_generic_type of CON_SCL_FCTR_D3_STATE : constant is 1;
    attribute mti_svvh_generic_type of PWR_DIS_D0_STATE : constant is 1;
    attribute mti_svvh_generic_type of DIS_SCL_FCTR_D0_STATE : constant is 1;
    attribute mti_svvh_generic_type of PWR_DIS_D1_STATE : constant is 1;
    attribute mti_svvh_generic_type of DIS_SCL_FCTR_D1_STATE : constant is 1;
    attribute mti_svvh_generic_type of PWR_DIS_D2_STATE : constant is 1;
    attribute mti_svvh_generic_type of DIS_SCL_FCTR_D2_STATE : constant is 1;
    attribute mti_svvh_generic_type of PWR_DIS_D3_STATE : constant is 1;
    attribute mti_svvh_generic_type of DIS_SCL_FCTR_D3_STATE : constant is 1;
    attribute mti_svvh_generic_type of CAL_BLK_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of SWAP_A_B_PAIRS : constant is 1;
    attribute mti_svvh_generic_type of INFINITECOMPLETIONS : constant is 1;
    attribute mti_svvh_generic_type of VC0_CREDITS_PH : constant is 1;
    attribute mti_svvh_generic_type of VC0_CREDITS_NPH : constant is 1;
    attribute mti_svvh_generic_type of CPL_STREAMING_PRIORITIZE_P_NP : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CLK : constant is 1;
    attribute mti_svvh_generic_type of TX_DIFF_BOOST : constant is 1;
    attribute mti_svvh_generic_type of TXDIFFCTRL : constant is 1;
    attribute mti_svvh_generic_type of TXBUFDIFFCTRL : constant is 1;
    attribute mti_svvh_generic_type of TXPREEMPHASIS : constant is 1;
    attribute mti_svvh_generic_type of GT_Debug_Ports : constant is 1;
    attribute mti_svvh_generic_type of GTDEBUGPORTS : constant is 1;
end endpoint_blk_plus_v1_15;
