library verilog;
use verilog.vl_types.all;
entity eth_mac_ram_sv_unit is
end eth_mac_ram_sv_unit;
